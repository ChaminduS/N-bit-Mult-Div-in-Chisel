module xor2(
  input   io_a,
  input   io_b,
  output  io_out
);
  assign io_out = io_a ^ io_b; // @[getOnesComplement.scala 13:20]
endmodule
module getOnesComplement(
  input         io_cin,
  input  [63:0] io_i1,
  output [63:0] io_onesComp
);
  wire  xor_0_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_0_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_0_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_1_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_1_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_1_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_2_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_2_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_2_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_3_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_3_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_3_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_4_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_4_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_4_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_5_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_5_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_5_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_6_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_6_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_6_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_7_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_7_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_7_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_8_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_8_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_8_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_9_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_9_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_9_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_10_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_10_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_10_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_11_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_11_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_11_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_12_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_12_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_12_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_13_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_13_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_13_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_14_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_14_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_14_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_15_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_15_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_15_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_16_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_16_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_16_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_17_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_17_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_17_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_18_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_18_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_18_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_19_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_19_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_19_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_20_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_20_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_20_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_21_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_21_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_21_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_22_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_22_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_22_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_23_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_23_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_23_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_24_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_24_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_24_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_25_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_25_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_25_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_26_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_26_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_26_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_27_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_27_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_27_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_28_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_28_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_28_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_29_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_29_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_29_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_30_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_30_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_30_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_31_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_31_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_31_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_32_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_32_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_32_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_33_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_33_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_33_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_34_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_34_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_34_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_35_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_35_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_35_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_36_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_36_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_36_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_37_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_37_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_37_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_38_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_38_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_38_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_39_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_39_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_39_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_40_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_40_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_40_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_41_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_41_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_41_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_42_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_42_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_42_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_43_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_43_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_43_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_44_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_44_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_44_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_45_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_45_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_45_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_46_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_46_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_46_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_47_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_47_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_47_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_48_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_48_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_48_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_49_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_49_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_49_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_50_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_50_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_50_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_51_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_51_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_51_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_52_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_52_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_52_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_53_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_53_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_53_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_54_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_54_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_54_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_55_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_55_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_55_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_56_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_56_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_56_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_57_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_57_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_57_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_58_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_58_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_58_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_59_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_59_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_59_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_60_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_60_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_60_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_61_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_61_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_61_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_62_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_62_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_62_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_63_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_63_io_b; // @[getOnesComplement.scala 24:33]
  wire  xor_63_io_out; // @[getOnesComplement.scala 24:33]
  wire [7:0] lo_lo_lo = {xor_7_io_out,xor_6_io_out,xor_5_io_out,xor_4_io_out,xor_3_io_out,xor_2_io_out,xor_1_io_out,
    xor_0_io_out}; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {xor_15_io_out,xor_14_io_out,xor_13_io_out,xor_12_io_out,xor_11_io_out,xor_10_io_out,xor_9_io_out,
    xor_8_io_out,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {xor_23_io_out,xor_22_io_out,xor_21_io_out,xor_20_io_out,xor_19_io_out,xor_18_io_out,
    xor_17_io_out,xor_16_io_out}; // @[Cat.scala 30:58]
  wire [31:0] lo = {xor_31_io_out,xor_30_io_out,xor_29_io_out,xor_28_io_out,xor_27_io_out,xor_26_io_out,xor_25_io_out,
    xor_24_io_out,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {xor_39_io_out,xor_38_io_out,xor_37_io_out,xor_36_io_out,xor_35_io_out,xor_34_io_out,
    xor_33_io_out,xor_32_io_out}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {xor_47_io_out,xor_46_io_out,xor_45_io_out,xor_44_io_out,xor_43_io_out,xor_42_io_out,xor_41_io_out
    ,xor_40_io_out,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {xor_55_io_out,xor_54_io_out,xor_53_io_out,xor_52_io_out,xor_51_io_out,xor_50_io_out,
    xor_49_io_out,xor_48_io_out}; // @[Cat.scala 30:58]
  wire [31:0] hi = {xor_63_io_out,xor_62_io_out,xor_61_io_out,xor_60_io_out,xor_59_io_out,xor_58_io_out,xor_57_io_out,
    xor_56_io_out,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  xor2 xor_0 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_0_io_a),
    .io_b(xor_0_io_b),
    .io_out(xor_0_io_out)
  );
  xor2 xor_1 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_1_io_a),
    .io_b(xor_1_io_b),
    .io_out(xor_1_io_out)
  );
  xor2 xor_2 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_2_io_a),
    .io_b(xor_2_io_b),
    .io_out(xor_2_io_out)
  );
  xor2 xor_3 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_3_io_a),
    .io_b(xor_3_io_b),
    .io_out(xor_3_io_out)
  );
  xor2 xor_4 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_4_io_a),
    .io_b(xor_4_io_b),
    .io_out(xor_4_io_out)
  );
  xor2 xor_5 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_5_io_a),
    .io_b(xor_5_io_b),
    .io_out(xor_5_io_out)
  );
  xor2 xor_6 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_6_io_a),
    .io_b(xor_6_io_b),
    .io_out(xor_6_io_out)
  );
  xor2 xor_7 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_7_io_a),
    .io_b(xor_7_io_b),
    .io_out(xor_7_io_out)
  );
  xor2 xor_8 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_8_io_a),
    .io_b(xor_8_io_b),
    .io_out(xor_8_io_out)
  );
  xor2 xor_9 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_9_io_a),
    .io_b(xor_9_io_b),
    .io_out(xor_9_io_out)
  );
  xor2 xor_10 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_10_io_a),
    .io_b(xor_10_io_b),
    .io_out(xor_10_io_out)
  );
  xor2 xor_11 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_11_io_a),
    .io_b(xor_11_io_b),
    .io_out(xor_11_io_out)
  );
  xor2 xor_12 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_12_io_a),
    .io_b(xor_12_io_b),
    .io_out(xor_12_io_out)
  );
  xor2 xor_13 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_13_io_a),
    .io_b(xor_13_io_b),
    .io_out(xor_13_io_out)
  );
  xor2 xor_14 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_14_io_a),
    .io_b(xor_14_io_b),
    .io_out(xor_14_io_out)
  );
  xor2 xor_15 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_15_io_a),
    .io_b(xor_15_io_b),
    .io_out(xor_15_io_out)
  );
  xor2 xor_16 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_16_io_a),
    .io_b(xor_16_io_b),
    .io_out(xor_16_io_out)
  );
  xor2 xor_17 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_17_io_a),
    .io_b(xor_17_io_b),
    .io_out(xor_17_io_out)
  );
  xor2 xor_18 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_18_io_a),
    .io_b(xor_18_io_b),
    .io_out(xor_18_io_out)
  );
  xor2 xor_19 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_19_io_a),
    .io_b(xor_19_io_b),
    .io_out(xor_19_io_out)
  );
  xor2 xor_20 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_20_io_a),
    .io_b(xor_20_io_b),
    .io_out(xor_20_io_out)
  );
  xor2 xor_21 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_21_io_a),
    .io_b(xor_21_io_b),
    .io_out(xor_21_io_out)
  );
  xor2 xor_22 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_22_io_a),
    .io_b(xor_22_io_b),
    .io_out(xor_22_io_out)
  );
  xor2 xor_23 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_23_io_a),
    .io_b(xor_23_io_b),
    .io_out(xor_23_io_out)
  );
  xor2 xor_24 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_24_io_a),
    .io_b(xor_24_io_b),
    .io_out(xor_24_io_out)
  );
  xor2 xor_25 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_25_io_a),
    .io_b(xor_25_io_b),
    .io_out(xor_25_io_out)
  );
  xor2 xor_26 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_26_io_a),
    .io_b(xor_26_io_b),
    .io_out(xor_26_io_out)
  );
  xor2 xor_27 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_27_io_a),
    .io_b(xor_27_io_b),
    .io_out(xor_27_io_out)
  );
  xor2 xor_28 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_28_io_a),
    .io_b(xor_28_io_b),
    .io_out(xor_28_io_out)
  );
  xor2 xor_29 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_29_io_a),
    .io_b(xor_29_io_b),
    .io_out(xor_29_io_out)
  );
  xor2 xor_30 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_30_io_a),
    .io_b(xor_30_io_b),
    .io_out(xor_30_io_out)
  );
  xor2 xor_31 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_31_io_a),
    .io_b(xor_31_io_b),
    .io_out(xor_31_io_out)
  );
  xor2 xor_32 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_32_io_a),
    .io_b(xor_32_io_b),
    .io_out(xor_32_io_out)
  );
  xor2 xor_33 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_33_io_a),
    .io_b(xor_33_io_b),
    .io_out(xor_33_io_out)
  );
  xor2 xor_34 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_34_io_a),
    .io_b(xor_34_io_b),
    .io_out(xor_34_io_out)
  );
  xor2 xor_35 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_35_io_a),
    .io_b(xor_35_io_b),
    .io_out(xor_35_io_out)
  );
  xor2 xor_36 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_36_io_a),
    .io_b(xor_36_io_b),
    .io_out(xor_36_io_out)
  );
  xor2 xor_37 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_37_io_a),
    .io_b(xor_37_io_b),
    .io_out(xor_37_io_out)
  );
  xor2 xor_38 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_38_io_a),
    .io_b(xor_38_io_b),
    .io_out(xor_38_io_out)
  );
  xor2 xor_39 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_39_io_a),
    .io_b(xor_39_io_b),
    .io_out(xor_39_io_out)
  );
  xor2 xor_40 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_40_io_a),
    .io_b(xor_40_io_b),
    .io_out(xor_40_io_out)
  );
  xor2 xor_41 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_41_io_a),
    .io_b(xor_41_io_b),
    .io_out(xor_41_io_out)
  );
  xor2 xor_42 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_42_io_a),
    .io_b(xor_42_io_b),
    .io_out(xor_42_io_out)
  );
  xor2 xor_43 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_43_io_a),
    .io_b(xor_43_io_b),
    .io_out(xor_43_io_out)
  );
  xor2 xor_44 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_44_io_a),
    .io_b(xor_44_io_b),
    .io_out(xor_44_io_out)
  );
  xor2 xor_45 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_45_io_a),
    .io_b(xor_45_io_b),
    .io_out(xor_45_io_out)
  );
  xor2 xor_46 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_46_io_a),
    .io_b(xor_46_io_b),
    .io_out(xor_46_io_out)
  );
  xor2 xor_47 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_47_io_a),
    .io_b(xor_47_io_b),
    .io_out(xor_47_io_out)
  );
  xor2 xor_48 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_48_io_a),
    .io_b(xor_48_io_b),
    .io_out(xor_48_io_out)
  );
  xor2 xor_49 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_49_io_a),
    .io_b(xor_49_io_b),
    .io_out(xor_49_io_out)
  );
  xor2 xor_50 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_50_io_a),
    .io_b(xor_50_io_b),
    .io_out(xor_50_io_out)
  );
  xor2 xor_51 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_51_io_a),
    .io_b(xor_51_io_b),
    .io_out(xor_51_io_out)
  );
  xor2 xor_52 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_52_io_a),
    .io_b(xor_52_io_b),
    .io_out(xor_52_io_out)
  );
  xor2 xor_53 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_53_io_a),
    .io_b(xor_53_io_b),
    .io_out(xor_53_io_out)
  );
  xor2 xor_54 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_54_io_a),
    .io_b(xor_54_io_b),
    .io_out(xor_54_io_out)
  );
  xor2 xor_55 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_55_io_a),
    .io_b(xor_55_io_b),
    .io_out(xor_55_io_out)
  );
  xor2 xor_56 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_56_io_a),
    .io_b(xor_56_io_b),
    .io_out(xor_56_io_out)
  );
  xor2 xor_57 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_57_io_a),
    .io_b(xor_57_io_b),
    .io_out(xor_57_io_out)
  );
  xor2 xor_58 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_58_io_a),
    .io_b(xor_58_io_b),
    .io_out(xor_58_io_out)
  );
  xor2 xor_59 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_59_io_a),
    .io_b(xor_59_io_b),
    .io_out(xor_59_io_out)
  );
  xor2 xor_60 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_60_io_a),
    .io_b(xor_60_io_b),
    .io_out(xor_60_io_out)
  );
  xor2 xor_61 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_61_io_a),
    .io_b(xor_61_io_b),
    .io_out(xor_61_io_out)
  );
  xor2 xor_62 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_62_io_a),
    .io_b(xor_62_io_b),
    .io_out(xor_62_io_out)
  );
  xor2 xor_63 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_63_io_a),
    .io_b(xor_63_io_b),
    .io_out(xor_63_io_out)
  );
  assign io_onesComp = {hi,lo}; // @[Cat.scala 30:58]
  assign xor_0_io_a = io_i1[0]; // @[getOnesComplement.scala 27:29]
  assign xor_0_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_1_io_a = io_i1[1]; // @[getOnesComplement.scala 27:29]
  assign xor_1_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_2_io_a = io_i1[2]; // @[getOnesComplement.scala 27:29]
  assign xor_2_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_3_io_a = io_i1[3]; // @[getOnesComplement.scala 27:29]
  assign xor_3_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_4_io_a = io_i1[4]; // @[getOnesComplement.scala 27:29]
  assign xor_4_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_5_io_a = io_i1[5]; // @[getOnesComplement.scala 27:29]
  assign xor_5_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_6_io_a = io_i1[6]; // @[getOnesComplement.scala 27:29]
  assign xor_6_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_7_io_a = io_i1[7]; // @[getOnesComplement.scala 27:29]
  assign xor_7_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_8_io_a = io_i1[8]; // @[getOnesComplement.scala 27:29]
  assign xor_8_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_9_io_a = io_i1[9]; // @[getOnesComplement.scala 27:29]
  assign xor_9_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_10_io_a = io_i1[10]; // @[getOnesComplement.scala 27:29]
  assign xor_10_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_11_io_a = io_i1[11]; // @[getOnesComplement.scala 27:29]
  assign xor_11_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_12_io_a = io_i1[12]; // @[getOnesComplement.scala 27:29]
  assign xor_12_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_13_io_a = io_i1[13]; // @[getOnesComplement.scala 27:29]
  assign xor_13_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_14_io_a = io_i1[14]; // @[getOnesComplement.scala 27:29]
  assign xor_14_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_15_io_a = io_i1[15]; // @[getOnesComplement.scala 27:29]
  assign xor_15_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_16_io_a = io_i1[16]; // @[getOnesComplement.scala 27:29]
  assign xor_16_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_17_io_a = io_i1[17]; // @[getOnesComplement.scala 27:29]
  assign xor_17_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_18_io_a = io_i1[18]; // @[getOnesComplement.scala 27:29]
  assign xor_18_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_19_io_a = io_i1[19]; // @[getOnesComplement.scala 27:29]
  assign xor_19_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_20_io_a = io_i1[20]; // @[getOnesComplement.scala 27:29]
  assign xor_20_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_21_io_a = io_i1[21]; // @[getOnesComplement.scala 27:29]
  assign xor_21_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_22_io_a = io_i1[22]; // @[getOnesComplement.scala 27:29]
  assign xor_22_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_23_io_a = io_i1[23]; // @[getOnesComplement.scala 27:29]
  assign xor_23_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_24_io_a = io_i1[24]; // @[getOnesComplement.scala 27:29]
  assign xor_24_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_25_io_a = io_i1[25]; // @[getOnesComplement.scala 27:29]
  assign xor_25_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_26_io_a = io_i1[26]; // @[getOnesComplement.scala 27:29]
  assign xor_26_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_27_io_a = io_i1[27]; // @[getOnesComplement.scala 27:29]
  assign xor_27_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_28_io_a = io_i1[28]; // @[getOnesComplement.scala 27:29]
  assign xor_28_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_29_io_a = io_i1[29]; // @[getOnesComplement.scala 27:29]
  assign xor_29_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_30_io_a = io_i1[30]; // @[getOnesComplement.scala 27:29]
  assign xor_30_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_31_io_a = io_i1[31]; // @[getOnesComplement.scala 27:29]
  assign xor_31_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_32_io_a = io_i1[32]; // @[getOnesComplement.scala 27:29]
  assign xor_32_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_33_io_a = io_i1[33]; // @[getOnesComplement.scala 27:29]
  assign xor_33_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_34_io_a = io_i1[34]; // @[getOnesComplement.scala 27:29]
  assign xor_34_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_35_io_a = io_i1[35]; // @[getOnesComplement.scala 27:29]
  assign xor_35_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_36_io_a = io_i1[36]; // @[getOnesComplement.scala 27:29]
  assign xor_36_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_37_io_a = io_i1[37]; // @[getOnesComplement.scala 27:29]
  assign xor_37_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_38_io_a = io_i1[38]; // @[getOnesComplement.scala 27:29]
  assign xor_38_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_39_io_a = io_i1[39]; // @[getOnesComplement.scala 27:29]
  assign xor_39_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_40_io_a = io_i1[40]; // @[getOnesComplement.scala 27:29]
  assign xor_40_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_41_io_a = io_i1[41]; // @[getOnesComplement.scala 27:29]
  assign xor_41_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_42_io_a = io_i1[42]; // @[getOnesComplement.scala 27:29]
  assign xor_42_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_43_io_a = io_i1[43]; // @[getOnesComplement.scala 27:29]
  assign xor_43_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_44_io_a = io_i1[44]; // @[getOnesComplement.scala 27:29]
  assign xor_44_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_45_io_a = io_i1[45]; // @[getOnesComplement.scala 27:29]
  assign xor_45_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_46_io_a = io_i1[46]; // @[getOnesComplement.scala 27:29]
  assign xor_46_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_47_io_a = io_i1[47]; // @[getOnesComplement.scala 27:29]
  assign xor_47_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_48_io_a = io_i1[48]; // @[getOnesComplement.scala 27:29]
  assign xor_48_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_49_io_a = io_i1[49]; // @[getOnesComplement.scala 27:29]
  assign xor_49_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_50_io_a = io_i1[50]; // @[getOnesComplement.scala 27:29]
  assign xor_50_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_51_io_a = io_i1[51]; // @[getOnesComplement.scala 27:29]
  assign xor_51_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_52_io_a = io_i1[52]; // @[getOnesComplement.scala 27:29]
  assign xor_52_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_53_io_a = io_i1[53]; // @[getOnesComplement.scala 27:29]
  assign xor_53_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_54_io_a = io_i1[54]; // @[getOnesComplement.scala 27:29]
  assign xor_54_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_55_io_a = io_i1[55]; // @[getOnesComplement.scala 27:29]
  assign xor_55_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_56_io_a = io_i1[56]; // @[getOnesComplement.scala 27:29]
  assign xor_56_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_57_io_a = io_i1[57]; // @[getOnesComplement.scala 27:29]
  assign xor_57_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_58_io_a = io_i1[58]; // @[getOnesComplement.scala 27:29]
  assign xor_58_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_59_io_a = io_i1[59]; // @[getOnesComplement.scala 27:29]
  assign xor_59_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_60_io_a = io_i1[60]; // @[getOnesComplement.scala 27:29]
  assign xor_60_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_61_io_a = io_i1[61]; // @[getOnesComplement.scala 27:29]
  assign xor_61_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_62_io_a = io_i1[62]; // @[getOnesComplement.scala 27:29]
  assign xor_62_io_b = io_cin; // @[getOnesComplement.scala 28:21]
  assign xor_63_io_a = io_i1[63]; // @[getOnesComplement.scala 27:29]
  assign xor_63_io_b = io_cin; // @[getOnesComplement.scala 28:21]
endmodule
module fullAdder(
  input   io_i0,
  input   io_i1,
  input   io_cin,
  output  io_sum,
  output  io_cout
);
  assign io_sum = io_i0 ^ io_i1 ^ io_cin; // @[addsub_64.scala 14:29]
  assign io_cout = io_i0 & io_i1 | io_i1 & io_cin | io_cin & io_i0; // @[addsub_64.scala 15:51]
endmodule
module addsub_64(
  input         io_cin,
  input  [63:0] io_onesComp_ip,
  input  [63:0] io_i0,
  output [63:0] io_sum
);
  wire  fa_0_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_0_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_0_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_0_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_0_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_1_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_1_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_1_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_1_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_1_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_2_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_2_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_2_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_2_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_2_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_3_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_3_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_3_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_3_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_3_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_4_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_4_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_4_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_4_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_4_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_5_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_5_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_5_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_5_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_5_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_6_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_6_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_6_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_6_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_6_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_7_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_7_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_7_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_7_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_7_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_8_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_8_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_8_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_8_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_8_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_9_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_9_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_9_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_9_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_9_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_10_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_10_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_10_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_10_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_10_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_11_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_11_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_11_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_11_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_11_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_12_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_12_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_12_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_12_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_12_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_13_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_13_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_13_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_13_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_13_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_14_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_14_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_14_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_14_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_14_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_15_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_15_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_15_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_15_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_15_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_16_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_16_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_16_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_16_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_16_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_17_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_17_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_17_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_17_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_17_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_18_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_18_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_18_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_18_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_18_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_19_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_19_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_19_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_19_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_19_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_20_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_20_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_20_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_20_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_20_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_21_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_21_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_21_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_21_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_21_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_22_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_22_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_22_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_22_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_22_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_23_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_23_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_23_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_23_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_23_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_24_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_24_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_24_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_24_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_24_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_25_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_25_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_25_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_25_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_25_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_26_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_26_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_26_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_26_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_26_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_27_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_27_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_27_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_27_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_27_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_28_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_28_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_28_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_28_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_28_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_29_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_29_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_29_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_29_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_29_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_30_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_30_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_30_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_30_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_30_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_31_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_31_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_31_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_31_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_31_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_32_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_32_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_32_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_32_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_32_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_33_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_33_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_33_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_33_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_33_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_34_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_34_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_34_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_34_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_34_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_35_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_35_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_35_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_35_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_35_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_36_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_36_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_36_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_36_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_36_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_37_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_37_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_37_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_37_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_37_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_38_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_38_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_38_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_38_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_38_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_39_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_39_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_39_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_39_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_39_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_40_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_40_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_40_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_40_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_40_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_41_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_41_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_41_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_41_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_41_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_42_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_42_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_42_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_42_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_42_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_43_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_43_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_43_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_43_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_43_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_44_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_44_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_44_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_44_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_44_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_45_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_45_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_45_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_45_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_45_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_46_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_46_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_46_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_46_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_46_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_47_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_47_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_47_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_47_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_47_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_48_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_48_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_48_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_48_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_48_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_49_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_49_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_49_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_49_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_49_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_50_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_50_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_50_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_50_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_50_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_51_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_51_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_51_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_51_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_51_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_52_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_52_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_52_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_52_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_52_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_53_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_53_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_53_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_53_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_53_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_54_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_54_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_54_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_54_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_54_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_55_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_55_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_55_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_55_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_55_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_56_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_56_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_56_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_56_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_56_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_57_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_57_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_57_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_57_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_57_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_58_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_58_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_58_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_58_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_58_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_59_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_59_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_59_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_59_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_59_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_60_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_60_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_60_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_60_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_60_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_61_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_61_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_61_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_61_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_61_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_62_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_62_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_62_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_62_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_62_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_63_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_63_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_63_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_63_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_63_io_cout; // @[addsub_64.scala 27:33]
  wire [7:0] lo_lo_lo = {fa_7_io_sum,fa_6_io_sum,fa_5_io_sum,fa_4_io_sum,fa_3_io_sum,fa_2_io_sum,fa_1_io_sum,fa_0_io_sum
    }; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {fa_15_io_sum,fa_14_io_sum,fa_13_io_sum,fa_12_io_sum,fa_11_io_sum,fa_10_io_sum,fa_9_io_sum,
    fa_8_io_sum,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {fa_23_io_sum,fa_22_io_sum,fa_21_io_sum,fa_20_io_sum,fa_19_io_sum,fa_18_io_sum,fa_17_io_sum,
    fa_16_io_sum}; // @[Cat.scala 30:58]
  wire [31:0] lo = {fa_31_io_sum,fa_30_io_sum,fa_29_io_sum,fa_28_io_sum,fa_27_io_sum,fa_26_io_sum,fa_25_io_sum,
    fa_24_io_sum,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {fa_39_io_sum,fa_38_io_sum,fa_37_io_sum,fa_36_io_sum,fa_35_io_sum,fa_34_io_sum,fa_33_io_sum,
    fa_32_io_sum}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {fa_47_io_sum,fa_46_io_sum,fa_45_io_sum,fa_44_io_sum,fa_43_io_sum,fa_42_io_sum,fa_41_io_sum,
    fa_40_io_sum,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {fa_55_io_sum,fa_54_io_sum,fa_53_io_sum,fa_52_io_sum,fa_51_io_sum,fa_50_io_sum,fa_49_io_sum,
    fa_48_io_sum}; // @[Cat.scala 30:58]
  wire [31:0] hi = {fa_63_io_sum,fa_62_io_sum,fa_61_io_sum,fa_60_io_sum,fa_59_io_sum,fa_58_io_sum,fa_57_io_sum,
    fa_56_io_sum,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  fullAdder fa_0 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_0_io_i0),
    .io_i1(fa_0_io_i1),
    .io_cin(fa_0_io_cin),
    .io_sum(fa_0_io_sum),
    .io_cout(fa_0_io_cout)
  );
  fullAdder fa_1 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_1_io_i0),
    .io_i1(fa_1_io_i1),
    .io_cin(fa_1_io_cin),
    .io_sum(fa_1_io_sum),
    .io_cout(fa_1_io_cout)
  );
  fullAdder fa_2 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_2_io_i0),
    .io_i1(fa_2_io_i1),
    .io_cin(fa_2_io_cin),
    .io_sum(fa_2_io_sum),
    .io_cout(fa_2_io_cout)
  );
  fullAdder fa_3 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_3_io_i0),
    .io_i1(fa_3_io_i1),
    .io_cin(fa_3_io_cin),
    .io_sum(fa_3_io_sum),
    .io_cout(fa_3_io_cout)
  );
  fullAdder fa_4 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_4_io_i0),
    .io_i1(fa_4_io_i1),
    .io_cin(fa_4_io_cin),
    .io_sum(fa_4_io_sum),
    .io_cout(fa_4_io_cout)
  );
  fullAdder fa_5 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_5_io_i0),
    .io_i1(fa_5_io_i1),
    .io_cin(fa_5_io_cin),
    .io_sum(fa_5_io_sum),
    .io_cout(fa_5_io_cout)
  );
  fullAdder fa_6 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_6_io_i0),
    .io_i1(fa_6_io_i1),
    .io_cin(fa_6_io_cin),
    .io_sum(fa_6_io_sum),
    .io_cout(fa_6_io_cout)
  );
  fullAdder fa_7 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_7_io_i0),
    .io_i1(fa_7_io_i1),
    .io_cin(fa_7_io_cin),
    .io_sum(fa_7_io_sum),
    .io_cout(fa_7_io_cout)
  );
  fullAdder fa_8 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_8_io_i0),
    .io_i1(fa_8_io_i1),
    .io_cin(fa_8_io_cin),
    .io_sum(fa_8_io_sum),
    .io_cout(fa_8_io_cout)
  );
  fullAdder fa_9 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_9_io_i0),
    .io_i1(fa_9_io_i1),
    .io_cin(fa_9_io_cin),
    .io_sum(fa_9_io_sum),
    .io_cout(fa_9_io_cout)
  );
  fullAdder fa_10 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_10_io_i0),
    .io_i1(fa_10_io_i1),
    .io_cin(fa_10_io_cin),
    .io_sum(fa_10_io_sum),
    .io_cout(fa_10_io_cout)
  );
  fullAdder fa_11 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_11_io_i0),
    .io_i1(fa_11_io_i1),
    .io_cin(fa_11_io_cin),
    .io_sum(fa_11_io_sum),
    .io_cout(fa_11_io_cout)
  );
  fullAdder fa_12 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_12_io_i0),
    .io_i1(fa_12_io_i1),
    .io_cin(fa_12_io_cin),
    .io_sum(fa_12_io_sum),
    .io_cout(fa_12_io_cout)
  );
  fullAdder fa_13 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_13_io_i0),
    .io_i1(fa_13_io_i1),
    .io_cin(fa_13_io_cin),
    .io_sum(fa_13_io_sum),
    .io_cout(fa_13_io_cout)
  );
  fullAdder fa_14 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_14_io_i0),
    .io_i1(fa_14_io_i1),
    .io_cin(fa_14_io_cin),
    .io_sum(fa_14_io_sum),
    .io_cout(fa_14_io_cout)
  );
  fullAdder fa_15 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_15_io_i0),
    .io_i1(fa_15_io_i1),
    .io_cin(fa_15_io_cin),
    .io_sum(fa_15_io_sum),
    .io_cout(fa_15_io_cout)
  );
  fullAdder fa_16 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_16_io_i0),
    .io_i1(fa_16_io_i1),
    .io_cin(fa_16_io_cin),
    .io_sum(fa_16_io_sum),
    .io_cout(fa_16_io_cout)
  );
  fullAdder fa_17 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_17_io_i0),
    .io_i1(fa_17_io_i1),
    .io_cin(fa_17_io_cin),
    .io_sum(fa_17_io_sum),
    .io_cout(fa_17_io_cout)
  );
  fullAdder fa_18 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_18_io_i0),
    .io_i1(fa_18_io_i1),
    .io_cin(fa_18_io_cin),
    .io_sum(fa_18_io_sum),
    .io_cout(fa_18_io_cout)
  );
  fullAdder fa_19 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_19_io_i0),
    .io_i1(fa_19_io_i1),
    .io_cin(fa_19_io_cin),
    .io_sum(fa_19_io_sum),
    .io_cout(fa_19_io_cout)
  );
  fullAdder fa_20 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_20_io_i0),
    .io_i1(fa_20_io_i1),
    .io_cin(fa_20_io_cin),
    .io_sum(fa_20_io_sum),
    .io_cout(fa_20_io_cout)
  );
  fullAdder fa_21 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_21_io_i0),
    .io_i1(fa_21_io_i1),
    .io_cin(fa_21_io_cin),
    .io_sum(fa_21_io_sum),
    .io_cout(fa_21_io_cout)
  );
  fullAdder fa_22 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_22_io_i0),
    .io_i1(fa_22_io_i1),
    .io_cin(fa_22_io_cin),
    .io_sum(fa_22_io_sum),
    .io_cout(fa_22_io_cout)
  );
  fullAdder fa_23 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_23_io_i0),
    .io_i1(fa_23_io_i1),
    .io_cin(fa_23_io_cin),
    .io_sum(fa_23_io_sum),
    .io_cout(fa_23_io_cout)
  );
  fullAdder fa_24 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_24_io_i0),
    .io_i1(fa_24_io_i1),
    .io_cin(fa_24_io_cin),
    .io_sum(fa_24_io_sum),
    .io_cout(fa_24_io_cout)
  );
  fullAdder fa_25 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_25_io_i0),
    .io_i1(fa_25_io_i1),
    .io_cin(fa_25_io_cin),
    .io_sum(fa_25_io_sum),
    .io_cout(fa_25_io_cout)
  );
  fullAdder fa_26 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_26_io_i0),
    .io_i1(fa_26_io_i1),
    .io_cin(fa_26_io_cin),
    .io_sum(fa_26_io_sum),
    .io_cout(fa_26_io_cout)
  );
  fullAdder fa_27 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_27_io_i0),
    .io_i1(fa_27_io_i1),
    .io_cin(fa_27_io_cin),
    .io_sum(fa_27_io_sum),
    .io_cout(fa_27_io_cout)
  );
  fullAdder fa_28 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_28_io_i0),
    .io_i1(fa_28_io_i1),
    .io_cin(fa_28_io_cin),
    .io_sum(fa_28_io_sum),
    .io_cout(fa_28_io_cout)
  );
  fullAdder fa_29 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_29_io_i0),
    .io_i1(fa_29_io_i1),
    .io_cin(fa_29_io_cin),
    .io_sum(fa_29_io_sum),
    .io_cout(fa_29_io_cout)
  );
  fullAdder fa_30 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_30_io_i0),
    .io_i1(fa_30_io_i1),
    .io_cin(fa_30_io_cin),
    .io_sum(fa_30_io_sum),
    .io_cout(fa_30_io_cout)
  );
  fullAdder fa_31 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_31_io_i0),
    .io_i1(fa_31_io_i1),
    .io_cin(fa_31_io_cin),
    .io_sum(fa_31_io_sum),
    .io_cout(fa_31_io_cout)
  );
  fullAdder fa_32 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_32_io_i0),
    .io_i1(fa_32_io_i1),
    .io_cin(fa_32_io_cin),
    .io_sum(fa_32_io_sum),
    .io_cout(fa_32_io_cout)
  );
  fullAdder fa_33 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_33_io_i0),
    .io_i1(fa_33_io_i1),
    .io_cin(fa_33_io_cin),
    .io_sum(fa_33_io_sum),
    .io_cout(fa_33_io_cout)
  );
  fullAdder fa_34 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_34_io_i0),
    .io_i1(fa_34_io_i1),
    .io_cin(fa_34_io_cin),
    .io_sum(fa_34_io_sum),
    .io_cout(fa_34_io_cout)
  );
  fullAdder fa_35 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_35_io_i0),
    .io_i1(fa_35_io_i1),
    .io_cin(fa_35_io_cin),
    .io_sum(fa_35_io_sum),
    .io_cout(fa_35_io_cout)
  );
  fullAdder fa_36 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_36_io_i0),
    .io_i1(fa_36_io_i1),
    .io_cin(fa_36_io_cin),
    .io_sum(fa_36_io_sum),
    .io_cout(fa_36_io_cout)
  );
  fullAdder fa_37 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_37_io_i0),
    .io_i1(fa_37_io_i1),
    .io_cin(fa_37_io_cin),
    .io_sum(fa_37_io_sum),
    .io_cout(fa_37_io_cout)
  );
  fullAdder fa_38 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_38_io_i0),
    .io_i1(fa_38_io_i1),
    .io_cin(fa_38_io_cin),
    .io_sum(fa_38_io_sum),
    .io_cout(fa_38_io_cout)
  );
  fullAdder fa_39 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_39_io_i0),
    .io_i1(fa_39_io_i1),
    .io_cin(fa_39_io_cin),
    .io_sum(fa_39_io_sum),
    .io_cout(fa_39_io_cout)
  );
  fullAdder fa_40 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_40_io_i0),
    .io_i1(fa_40_io_i1),
    .io_cin(fa_40_io_cin),
    .io_sum(fa_40_io_sum),
    .io_cout(fa_40_io_cout)
  );
  fullAdder fa_41 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_41_io_i0),
    .io_i1(fa_41_io_i1),
    .io_cin(fa_41_io_cin),
    .io_sum(fa_41_io_sum),
    .io_cout(fa_41_io_cout)
  );
  fullAdder fa_42 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_42_io_i0),
    .io_i1(fa_42_io_i1),
    .io_cin(fa_42_io_cin),
    .io_sum(fa_42_io_sum),
    .io_cout(fa_42_io_cout)
  );
  fullAdder fa_43 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_43_io_i0),
    .io_i1(fa_43_io_i1),
    .io_cin(fa_43_io_cin),
    .io_sum(fa_43_io_sum),
    .io_cout(fa_43_io_cout)
  );
  fullAdder fa_44 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_44_io_i0),
    .io_i1(fa_44_io_i1),
    .io_cin(fa_44_io_cin),
    .io_sum(fa_44_io_sum),
    .io_cout(fa_44_io_cout)
  );
  fullAdder fa_45 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_45_io_i0),
    .io_i1(fa_45_io_i1),
    .io_cin(fa_45_io_cin),
    .io_sum(fa_45_io_sum),
    .io_cout(fa_45_io_cout)
  );
  fullAdder fa_46 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_46_io_i0),
    .io_i1(fa_46_io_i1),
    .io_cin(fa_46_io_cin),
    .io_sum(fa_46_io_sum),
    .io_cout(fa_46_io_cout)
  );
  fullAdder fa_47 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_47_io_i0),
    .io_i1(fa_47_io_i1),
    .io_cin(fa_47_io_cin),
    .io_sum(fa_47_io_sum),
    .io_cout(fa_47_io_cout)
  );
  fullAdder fa_48 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_48_io_i0),
    .io_i1(fa_48_io_i1),
    .io_cin(fa_48_io_cin),
    .io_sum(fa_48_io_sum),
    .io_cout(fa_48_io_cout)
  );
  fullAdder fa_49 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_49_io_i0),
    .io_i1(fa_49_io_i1),
    .io_cin(fa_49_io_cin),
    .io_sum(fa_49_io_sum),
    .io_cout(fa_49_io_cout)
  );
  fullAdder fa_50 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_50_io_i0),
    .io_i1(fa_50_io_i1),
    .io_cin(fa_50_io_cin),
    .io_sum(fa_50_io_sum),
    .io_cout(fa_50_io_cout)
  );
  fullAdder fa_51 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_51_io_i0),
    .io_i1(fa_51_io_i1),
    .io_cin(fa_51_io_cin),
    .io_sum(fa_51_io_sum),
    .io_cout(fa_51_io_cout)
  );
  fullAdder fa_52 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_52_io_i0),
    .io_i1(fa_52_io_i1),
    .io_cin(fa_52_io_cin),
    .io_sum(fa_52_io_sum),
    .io_cout(fa_52_io_cout)
  );
  fullAdder fa_53 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_53_io_i0),
    .io_i1(fa_53_io_i1),
    .io_cin(fa_53_io_cin),
    .io_sum(fa_53_io_sum),
    .io_cout(fa_53_io_cout)
  );
  fullAdder fa_54 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_54_io_i0),
    .io_i1(fa_54_io_i1),
    .io_cin(fa_54_io_cin),
    .io_sum(fa_54_io_sum),
    .io_cout(fa_54_io_cout)
  );
  fullAdder fa_55 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_55_io_i0),
    .io_i1(fa_55_io_i1),
    .io_cin(fa_55_io_cin),
    .io_sum(fa_55_io_sum),
    .io_cout(fa_55_io_cout)
  );
  fullAdder fa_56 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_56_io_i0),
    .io_i1(fa_56_io_i1),
    .io_cin(fa_56_io_cin),
    .io_sum(fa_56_io_sum),
    .io_cout(fa_56_io_cout)
  );
  fullAdder fa_57 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_57_io_i0),
    .io_i1(fa_57_io_i1),
    .io_cin(fa_57_io_cin),
    .io_sum(fa_57_io_sum),
    .io_cout(fa_57_io_cout)
  );
  fullAdder fa_58 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_58_io_i0),
    .io_i1(fa_58_io_i1),
    .io_cin(fa_58_io_cin),
    .io_sum(fa_58_io_sum),
    .io_cout(fa_58_io_cout)
  );
  fullAdder fa_59 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_59_io_i0),
    .io_i1(fa_59_io_i1),
    .io_cin(fa_59_io_cin),
    .io_sum(fa_59_io_sum),
    .io_cout(fa_59_io_cout)
  );
  fullAdder fa_60 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_60_io_i0),
    .io_i1(fa_60_io_i1),
    .io_cin(fa_60_io_cin),
    .io_sum(fa_60_io_sum),
    .io_cout(fa_60_io_cout)
  );
  fullAdder fa_61 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_61_io_i0),
    .io_i1(fa_61_io_i1),
    .io_cin(fa_61_io_cin),
    .io_sum(fa_61_io_sum),
    .io_cout(fa_61_io_cout)
  );
  fullAdder fa_62 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_62_io_i0),
    .io_i1(fa_62_io_i1),
    .io_cin(fa_62_io_cin),
    .io_sum(fa_62_io_sum),
    .io_cout(fa_62_io_cout)
  );
  fullAdder fa_63 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_63_io_i0),
    .io_i1(fa_63_io_i1),
    .io_cin(fa_63_io_cin),
    .io_sum(fa_63_io_sum),
    .io_cout(fa_63_io_cout)
  );
  assign io_sum = {hi,lo}; // @[Cat.scala 30:58]
  assign fa_0_io_i0 = io_i0[0]; // @[addsub_64.scala 30:25]
  assign fa_0_io_i1 = io_onesComp_ip[0]; // @[addsub_64.scala 31:34]
  assign fa_0_io_cin = io_cin; // @[addsub_64.scala 32:18]
  assign fa_1_io_i0 = io_i0[1]; // @[addsub_64.scala 36:29]
  assign fa_1_io_i1 = io_onesComp_ip[1]; // @[addsub_64.scala 37:38]
  assign fa_1_io_cin = fa_0_io_cout; // @[addsub_64.scala 38:22]
  assign fa_2_io_i0 = io_i0[2]; // @[addsub_64.scala 36:29]
  assign fa_2_io_i1 = io_onesComp_ip[2]; // @[addsub_64.scala 37:38]
  assign fa_2_io_cin = fa_1_io_cout; // @[addsub_64.scala 38:22]
  assign fa_3_io_i0 = io_i0[3]; // @[addsub_64.scala 36:29]
  assign fa_3_io_i1 = io_onesComp_ip[3]; // @[addsub_64.scala 37:38]
  assign fa_3_io_cin = fa_2_io_cout; // @[addsub_64.scala 38:22]
  assign fa_4_io_i0 = io_i0[4]; // @[addsub_64.scala 36:29]
  assign fa_4_io_i1 = io_onesComp_ip[4]; // @[addsub_64.scala 37:38]
  assign fa_4_io_cin = fa_3_io_cout; // @[addsub_64.scala 38:22]
  assign fa_5_io_i0 = io_i0[5]; // @[addsub_64.scala 36:29]
  assign fa_5_io_i1 = io_onesComp_ip[5]; // @[addsub_64.scala 37:38]
  assign fa_5_io_cin = fa_4_io_cout; // @[addsub_64.scala 38:22]
  assign fa_6_io_i0 = io_i0[6]; // @[addsub_64.scala 36:29]
  assign fa_6_io_i1 = io_onesComp_ip[6]; // @[addsub_64.scala 37:38]
  assign fa_6_io_cin = fa_5_io_cout; // @[addsub_64.scala 38:22]
  assign fa_7_io_i0 = io_i0[7]; // @[addsub_64.scala 36:29]
  assign fa_7_io_i1 = io_onesComp_ip[7]; // @[addsub_64.scala 37:38]
  assign fa_7_io_cin = fa_6_io_cout; // @[addsub_64.scala 38:22]
  assign fa_8_io_i0 = io_i0[8]; // @[addsub_64.scala 36:29]
  assign fa_8_io_i1 = io_onesComp_ip[8]; // @[addsub_64.scala 37:38]
  assign fa_8_io_cin = fa_7_io_cout; // @[addsub_64.scala 38:22]
  assign fa_9_io_i0 = io_i0[9]; // @[addsub_64.scala 36:29]
  assign fa_9_io_i1 = io_onesComp_ip[9]; // @[addsub_64.scala 37:38]
  assign fa_9_io_cin = fa_8_io_cout; // @[addsub_64.scala 38:22]
  assign fa_10_io_i0 = io_i0[10]; // @[addsub_64.scala 36:29]
  assign fa_10_io_i1 = io_onesComp_ip[10]; // @[addsub_64.scala 37:38]
  assign fa_10_io_cin = fa_9_io_cout; // @[addsub_64.scala 38:22]
  assign fa_11_io_i0 = io_i0[11]; // @[addsub_64.scala 36:29]
  assign fa_11_io_i1 = io_onesComp_ip[11]; // @[addsub_64.scala 37:38]
  assign fa_11_io_cin = fa_10_io_cout; // @[addsub_64.scala 38:22]
  assign fa_12_io_i0 = io_i0[12]; // @[addsub_64.scala 36:29]
  assign fa_12_io_i1 = io_onesComp_ip[12]; // @[addsub_64.scala 37:38]
  assign fa_12_io_cin = fa_11_io_cout; // @[addsub_64.scala 38:22]
  assign fa_13_io_i0 = io_i0[13]; // @[addsub_64.scala 36:29]
  assign fa_13_io_i1 = io_onesComp_ip[13]; // @[addsub_64.scala 37:38]
  assign fa_13_io_cin = fa_12_io_cout; // @[addsub_64.scala 38:22]
  assign fa_14_io_i0 = io_i0[14]; // @[addsub_64.scala 36:29]
  assign fa_14_io_i1 = io_onesComp_ip[14]; // @[addsub_64.scala 37:38]
  assign fa_14_io_cin = fa_13_io_cout; // @[addsub_64.scala 38:22]
  assign fa_15_io_i0 = io_i0[15]; // @[addsub_64.scala 36:29]
  assign fa_15_io_i1 = io_onesComp_ip[15]; // @[addsub_64.scala 37:38]
  assign fa_15_io_cin = fa_14_io_cout; // @[addsub_64.scala 38:22]
  assign fa_16_io_i0 = io_i0[16]; // @[addsub_64.scala 36:29]
  assign fa_16_io_i1 = io_onesComp_ip[16]; // @[addsub_64.scala 37:38]
  assign fa_16_io_cin = fa_15_io_cout; // @[addsub_64.scala 38:22]
  assign fa_17_io_i0 = io_i0[17]; // @[addsub_64.scala 36:29]
  assign fa_17_io_i1 = io_onesComp_ip[17]; // @[addsub_64.scala 37:38]
  assign fa_17_io_cin = fa_16_io_cout; // @[addsub_64.scala 38:22]
  assign fa_18_io_i0 = io_i0[18]; // @[addsub_64.scala 36:29]
  assign fa_18_io_i1 = io_onesComp_ip[18]; // @[addsub_64.scala 37:38]
  assign fa_18_io_cin = fa_17_io_cout; // @[addsub_64.scala 38:22]
  assign fa_19_io_i0 = io_i0[19]; // @[addsub_64.scala 36:29]
  assign fa_19_io_i1 = io_onesComp_ip[19]; // @[addsub_64.scala 37:38]
  assign fa_19_io_cin = fa_18_io_cout; // @[addsub_64.scala 38:22]
  assign fa_20_io_i0 = io_i0[20]; // @[addsub_64.scala 36:29]
  assign fa_20_io_i1 = io_onesComp_ip[20]; // @[addsub_64.scala 37:38]
  assign fa_20_io_cin = fa_19_io_cout; // @[addsub_64.scala 38:22]
  assign fa_21_io_i0 = io_i0[21]; // @[addsub_64.scala 36:29]
  assign fa_21_io_i1 = io_onesComp_ip[21]; // @[addsub_64.scala 37:38]
  assign fa_21_io_cin = fa_20_io_cout; // @[addsub_64.scala 38:22]
  assign fa_22_io_i0 = io_i0[22]; // @[addsub_64.scala 36:29]
  assign fa_22_io_i1 = io_onesComp_ip[22]; // @[addsub_64.scala 37:38]
  assign fa_22_io_cin = fa_21_io_cout; // @[addsub_64.scala 38:22]
  assign fa_23_io_i0 = io_i0[23]; // @[addsub_64.scala 36:29]
  assign fa_23_io_i1 = io_onesComp_ip[23]; // @[addsub_64.scala 37:38]
  assign fa_23_io_cin = fa_22_io_cout; // @[addsub_64.scala 38:22]
  assign fa_24_io_i0 = io_i0[24]; // @[addsub_64.scala 36:29]
  assign fa_24_io_i1 = io_onesComp_ip[24]; // @[addsub_64.scala 37:38]
  assign fa_24_io_cin = fa_23_io_cout; // @[addsub_64.scala 38:22]
  assign fa_25_io_i0 = io_i0[25]; // @[addsub_64.scala 36:29]
  assign fa_25_io_i1 = io_onesComp_ip[25]; // @[addsub_64.scala 37:38]
  assign fa_25_io_cin = fa_24_io_cout; // @[addsub_64.scala 38:22]
  assign fa_26_io_i0 = io_i0[26]; // @[addsub_64.scala 36:29]
  assign fa_26_io_i1 = io_onesComp_ip[26]; // @[addsub_64.scala 37:38]
  assign fa_26_io_cin = fa_25_io_cout; // @[addsub_64.scala 38:22]
  assign fa_27_io_i0 = io_i0[27]; // @[addsub_64.scala 36:29]
  assign fa_27_io_i1 = io_onesComp_ip[27]; // @[addsub_64.scala 37:38]
  assign fa_27_io_cin = fa_26_io_cout; // @[addsub_64.scala 38:22]
  assign fa_28_io_i0 = io_i0[28]; // @[addsub_64.scala 36:29]
  assign fa_28_io_i1 = io_onesComp_ip[28]; // @[addsub_64.scala 37:38]
  assign fa_28_io_cin = fa_27_io_cout; // @[addsub_64.scala 38:22]
  assign fa_29_io_i0 = io_i0[29]; // @[addsub_64.scala 36:29]
  assign fa_29_io_i1 = io_onesComp_ip[29]; // @[addsub_64.scala 37:38]
  assign fa_29_io_cin = fa_28_io_cout; // @[addsub_64.scala 38:22]
  assign fa_30_io_i0 = io_i0[30]; // @[addsub_64.scala 36:29]
  assign fa_30_io_i1 = io_onesComp_ip[30]; // @[addsub_64.scala 37:38]
  assign fa_30_io_cin = fa_29_io_cout; // @[addsub_64.scala 38:22]
  assign fa_31_io_i0 = io_i0[31]; // @[addsub_64.scala 36:29]
  assign fa_31_io_i1 = io_onesComp_ip[31]; // @[addsub_64.scala 37:38]
  assign fa_31_io_cin = fa_30_io_cout; // @[addsub_64.scala 38:22]
  assign fa_32_io_i0 = io_i0[32]; // @[addsub_64.scala 36:29]
  assign fa_32_io_i1 = io_onesComp_ip[32]; // @[addsub_64.scala 37:38]
  assign fa_32_io_cin = fa_31_io_cout; // @[addsub_64.scala 38:22]
  assign fa_33_io_i0 = io_i0[33]; // @[addsub_64.scala 36:29]
  assign fa_33_io_i1 = io_onesComp_ip[33]; // @[addsub_64.scala 37:38]
  assign fa_33_io_cin = fa_32_io_cout; // @[addsub_64.scala 38:22]
  assign fa_34_io_i0 = io_i0[34]; // @[addsub_64.scala 36:29]
  assign fa_34_io_i1 = io_onesComp_ip[34]; // @[addsub_64.scala 37:38]
  assign fa_34_io_cin = fa_33_io_cout; // @[addsub_64.scala 38:22]
  assign fa_35_io_i0 = io_i0[35]; // @[addsub_64.scala 36:29]
  assign fa_35_io_i1 = io_onesComp_ip[35]; // @[addsub_64.scala 37:38]
  assign fa_35_io_cin = fa_34_io_cout; // @[addsub_64.scala 38:22]
  assign fa_36_io_i0 = io_i0[36]; // @[addsub_64.scala 36:29]
  assign fa_36_io_i1 = io_onesComp_ip[36]; // @[addsub_64.scala 37:38]
  assign fa_36_io_cin = fa_35_io_cout; // @[addsub_64.scala 38:22]
  assign fa_37_io_i0 = io_i0[37]; // @[addsub_64.scala 36:29]
  assign fa_37_io_i1 = io_onesComp_ip[37]; // @[addsub_64.scala 37:38]
  assign fa_37_io_cin = fa_36_io_cout; // @[addsub_64.scala 38:22]
  assign fa_38_io_i0 = io_i0[38]; // @[addsub_64.scala 36:29]
  assign fa_38_io_i1 = io_onesComp_ip[38]; // @[addsub_64.scala 37:38]
  assign fa_38_io_cin = fa_37_io_cout; // @[addsub_64.scala 38:22]
  assign fa_39_io_i0 = io_i0[39]; // @[addsub_64.scala 36:29]
  assign fa_39_io_i1 = io_onesComp_ip[39]; // @[addsub_64.scala 37:38]
  assign fa_39_io_cin = fa_38_io_cout; // @[addsub_64.scala 38:22]
  assign fa_40_io_i0 = io_i0[40]; // @[addsub_64.scala 36:29]
  assign fa_40_io_i1 = io_onesComp_ip[40]; // @[addsub_64.scala 37:38]
  assign fa_40_io_cin = fa_39_io_cout; // @[addsub_64.scala 38:22]
  assign fa_41_io_i0 = io_i0[41]; // @[addsub_64.scala 36:29]
  assign fa_41_io_i1 = io_onesComp_ip[41]; // @[addsub_64.scala 37:38]
  assign fa_41_io_cin = fa_40_io_cout; // @[addsub_64.scala 38:22]
  assign fa_42_io_i0 = io_i0[42]; // @[addsub_64.scala 36:29]
  assign fa_42_io_i1 = io_onesComp_ip[42]; // @[addsub_64.scala 37:38]
  assign fa_42_io_cin = fa_41_io_cout; // @[addsub_64.scala 38:22]
  assign fa_43_io_i0 = io_i0[43]; // @[addsub_64.scala 36:29]
  assign fa_43_io_i1 = io_onesComp_ip[43]; // @[addsub_64.scala 37:38]
  assign fa_43_io_cin = fa_42_io_cout; // @[addsub_64.scala 38:22]
  assign fa_44_io_i0 = io_i0[44]; // @[addsub_64.scala 36:29]
  assign fa_44_io_i1 = io_onesComp_ip[44]; // @[addsub_64.scala 37:38]
  assign fa_44_io_cin = fa_43_io_cout; // @[addsub_64.scala 38:22]
  assign fa_45_io_i0 = io_i0[45]; // @[addsub_64.scala 36:29]
  assign fa_45_io_i1 = io_onesComp_ip[45]; // @[addsub_64.scala 37:38]
  assign fa_45_io_cin = fa_44_io_cout; // @[addsub_64.scala 38:22]
  assign fa_46_io_i0 = io_i0[46]; // @[addsub_64.scala 36:29]
  assign fa_46_io_i1 = io_onesComp_ip[46]; // @[addsub_64.scala 37:38]
  assign fa_46_io_cin = fa_45_io_cout; // @[addsub_64.scala 38:22]
  assign fa_47_io_i0 = io_i0[47]; // @[addsub_64.scala 36:29]
  assign fa_47_io_i1 = io_onesComp_ip[47]; // @[addsub_64.scala 37:38]
  assign fa_47_io_cin = fa_46_io_cout; // @[addsub_64.scala 38:22]
  assign fa_48_io_i0 = io_i0[48]; // @[addsub_64.scala 36:29]
  assign fa_48_io_i1 = io_onesComp_ip[48]; // @[addsub_64.scala 37:38]
  assign fa_48_io_cin = fa_47_io_cout; // @[addsub_64.scala 38:22]
  assign fa_49_io_i0 = io_i0[49]; // @[addsub_64.scala 36:29]
  assign fa_49_io_i1 = io_onesComp_ip[49]; // @[addsub_64.scala 37:38]
  assign fa_49_io_cin = fa_48_io_cout; // @[addsub_64.scala 38:22]
  assign fa_50_io_i0 = io_i0[50]; // @[addsub_64.scala 36:29]
  assign fa_50_io_i1 = io_onesComp_ip[50]; // @[addsub_64.scala 37:38]
  assign fa_50_io_cin = fa_49_io_cout; // @[addsub_64.scala 38:22]
  assign fa_51_io_i0 = io_i0[51]; // @[addsub_64.scala 36:29]
  assign fa_51_io_i1 = io_onesComp_ip[51]; // @[addsub_64.scala 37:38]
  assign fa_51_io_cin = fa_50_io_cout; // @[addsub_64.scala 38:22]
  assign fa_52_io_i0 = io_i0[52]; // @[addsub_64.scala 36:29]
  assign fa_52_io_i1 = io_onesComp_ip[52]; // @[addsub_64.scala 37:38]
  assign fa_52_io_cin = fa_51_io_cout; // @[addsub_64.scala 38:22]
  assign fa_53_io_i0 = io_i0[53]; // @[addsub_64.scala 36:29]
  assign fa_53_io_i1 = io_onesComp_ip[53]; // @[addsub_64.scala 37:38]
  assign fa_53_io_cin = fa_52_io_cout; // @[addsub_64.scala 38:22]
  assign fa_54_io_i0 = io_i0[54]; // @[addsub_64.scala 36:29]
  assign fa_54_io_i1 = io_onesComp_ip[54]; // @[addsub_64.scala 37:38]
  assign fa_54_io_cin = fa_53_io_cout; // @[addsub_64.scala 38:22]
  assign fa_55_io_i0 = io_i0[55]; // @[addsub_64.scala 36:29]
  assign fa_55_io_i1 = io_onesComp_ip[55]; // @[addsub_64.scala 37:38]
  assign fa_55_io_cin = fa_54_io_cout; // @[addsub_64.scala 38:22]
  assign fa_56_io_i0 = io_i0[56]; // @[addsub_64.scala 36:29]
  assign fa_56_io_i1 = io_onesComp_ip[56]; // @[addsub_64.scala 37:38]
  assign fa_56_io_cin = fa_55_io_cout; // @[addsub_64.scala 38:22]
  assign fa_57_io_i0 = io_i0[57]; // @[addsub_64.scala 36:29]
  assign fa_57_io_i1 = io_onesComp_ip[57]; // @[addsub_64.scala 37:38]
  assign fa_57_io_cin = fa_56_io_cout; // @[addsub_64.scala 38:22]
  assign fa_58_io_i0 = io_i0[58]; // @[addsub_64.scala 36:29]
  assign fa_58_io_i1 = io_onesComp_ip[58]; // @[addsub_64.scala 37:38]
  assign fa_58_io_cin = fa_57_io_cout; // @[addsub_64.scala 38:22]
  assign fa_59_io_i0 = io_i0[59]; // @[addsub_64.scala 36:29]
  assign fa_59_io_i1 = io_onesComp_ip[59]; // @[addsub_64.scala 37:38]
  assign fa_59_io_cin = fa_58_io_cout; // @[addsub_64.scala 38:22]
  assign fa_60_io_i0 = io_i0[60]; // @[addsub_64.scala 36:29]
  assign fa_60_io_i1 = io_onesComp_ip[60]; // @[addsub_64.scala 37:38]
  assign fa_60_io_cin = fa_59_io_cout; // @[addsub_64.scala 38:22]
  assign fa_61_io_i0 = io_i0[61]; // @[addsub_64.scala 36:29]
  assign fa_61_io_i1 = io_onesComp_ip[61]; // @[addsub_64.scala 37:38]
  assign fa_61_io_cin = fa_60_io_cout; // @[addsub_64.scala 38:22]
  assign fa_62_io_i0 = io_i0[62]; // @[addsub_64.scala 36:29]
  assign fa_62_io_i1 = io_onesComp_ip[62]; // @[addsub_64.scala 37:38]
  assign fa_62_io_cin = fa_61_io_cout; // @[addsub_64.scala 38:22]
  assign fa_63_io_i0 = io_i0[63]; // @[addsub_64.scala 36:29]
  assign fa_63_io_i1 = io_onesComp_ip[63]; // @[addsub_64.scala 37:38]
  assign fa_63_io_cin = fa_62_io_cout; // @[addsub_64.scala 38:22]
endmodule
module booth_substep(
  input  [63:0] io_acc,
  input  [63:0] io_Q,
  input         io_q0,
  input  [63:0] io_multiplicand,
  output [63:0] io_next_acc,
  output [63:0] io_next_Q,
  output        io_q0_next
);
  wire  g0_io_cin; // @[booth_substep.scala 17:20]
  wire [63:0] g0_io_i1; // @[booth_substep.scala 17:20]
  wire [63:0] g0_io_onesComp; // @[booth_substep.scala 17:20]
  wire  as0_io_cin; // @[booth_substep.scala 27:21]
  wire [63:0] as0_io_onesComp_ip; // @[booth_substep.scala 27:21]
  wire [63:0] as0_io_i0; // @[booth_substep.scala 27:21]
  wire [63:0] as0_io_sum; // @[booth_substep.scala 27:21]
  wire [63:0] _T_3 = io_acc; // @[booth_substep.scala 33:25]
  wire [63:0] _T_7 = io_Q; // @[booth_substep.scala 46:29]
  wire [63:0] addsub_temp = as0_io_sum; // @[booth_substep.scala 29:27 booth_substep.scala 34:17]
  wire [62:0] next_Q_temp = io_Q[0] == io_q0 ? _T_7[63:1] : _T_7[63:1]; // @[booth_substep.scala 44:29 booth_substep.scala 46:21 booth_substep.scala 56:21]
  wire  next_Q_MSB = io_Q[0] == io_q0 ? io_acc[0] : addsub_temp[0]; // @[booth_substep.scala 44:29 booth_substep.scala 47:20 booth_substep.scala 57:20]
  wire [62:0] next_acc_temp = io_Q[0] == io_q0 ? _T_3[63:1] : addsub_temp[63:1]; // @[booth_substep.scala 44:29 booth_substep.scala 48:23 booth_substep.scala 58:23]
  wire  next_acc_MSB = io_Q[0] == io_q0 ? io_acc[63] : addsub_temp[63]; // @[booth_substep.scala 44:29]
  getOnesComplement g0 ( // @[booth_substep.scala 17:20]
    .io_cin(g0_io_cin),
    .io_i1(g0_io_i1),
    .io_onesComp(g0_io_onesComp)
  );
  addsub_64 as0 ( // @[booth_substep.scala 27:21]
    .io_cin(as0_io_cin),
    .io_onesComp_ip(as0_io_onesComp_ip),
    .io_i0(as0_io_i0),
    .io_sum(as0_io_sum)
  );
  assign io_next_acc = {next_acc_MSB,next_acc_temp}; // @[booth_substep.scala 67:53]
  assign io_next_Q = {next_Q_MSB,next_Q_temp}; // @[booth_substep.scala 66:47]
  assign io_q0_next = io_Q[0] == io_q0 ? io_Q[0] : io_Q[0]; // @[booth_substep.scala 44:29 booth_substep.scala 45:20 booth_substep.scala 55:20]
  assign g0_io_cin = io_Q[0]; // @[booth_substep.scala 21:22]
  assign g0_io_i1 = io_multiplicand; // @[booth_substep.scala 22:33]
  assign as0_io_cin = io_Q[0]; // @[booth_substep.scala 31:23]
  assign as0_io_onesComp_ip = g0_io_onesComp; // @[booth_substep.scala 19:22 booth_substep.scala 23:12]
  assign as0_io_i0 = io_acc; // @[booth_substep.scala 33:25]
endmodule
module booth_multiplier(
  input          clock,
  input          reset,
  input  [63:0]  io_multiplier,
  input  [63:0]  io_multiplicand,
  output [127:0] io_product
);
  wire [63:0] bs_0_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_0_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_0_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_0_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_0_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_0_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_0_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_1_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_1_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_1_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_1_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_1_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_1_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_1_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_2_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_2_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_2_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_2_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_2_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_2_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_2_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_3_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_3_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_3_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_3_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_3_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_3_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_3_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_4_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_4_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_4_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_4_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_4_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_4_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_4_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_5_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_5_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_5_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_5_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_5_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_5_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_5_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_6_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_6_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_6_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_6_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_6_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_6_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_6_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_7_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_7_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_7_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_7_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_7_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_7_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_7_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_8_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_8_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_8_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_8_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_8_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_8_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_8_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_9_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_9_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_9_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_9_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_9_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_9_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_9_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_10_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_10_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_10_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_10_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_10_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_10_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_10_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_11_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_11_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_11_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_11_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_11_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_11_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_11_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_12_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_12_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_12_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_12_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_12_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_12_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_12_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_13_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_13_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_13_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_13_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_13_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_13_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_13_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_14_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_14_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_14_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_14_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_14_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_14_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_14_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_15_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_15_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_15_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_15_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_15_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_15_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_15_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_16_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_16_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_16_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_16_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_16_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_16_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_16_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_17_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_17_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_17_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_17_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_17_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_17_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_17_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_18_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_18_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_18_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_18_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_18_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_18_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_18_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_19_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_19_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_19_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_19_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_19_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_19_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_19_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_20_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_20_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_20_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_20_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_20_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_20_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_20_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_21_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_21_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_21_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_21_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_21_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_21_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_21_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_22_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_22_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_22_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_22_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_22_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_22_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_22_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_23_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_23_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_23_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_23_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_23_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_23_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_23_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_24_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_24_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_24_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_24_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_24_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_24_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_24_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_25_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_25_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_25_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_25_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_25_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_25_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_25_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_26_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_26_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_26_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_26_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_26_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_26_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_26_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_27_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_27_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_27_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_27_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_27_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_27_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_27_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_28_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_28_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_28_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_28_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_28_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_28_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_28_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_29_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_29_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_29_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_29_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_29_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_29_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_29_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_30_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_30_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_30_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_30_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_30_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_30_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_30_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_31_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_31_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_31_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_31_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_31_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_31_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_31_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_32_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_32_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_32_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_32_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_32_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_32_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_32_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_33_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_33_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_33_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_33_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_33_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_33_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_33_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_34_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_34_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_34_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_34_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_34_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_34_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_34_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_35_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_35_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_35_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_35_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_35_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_35_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_35_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_36_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_36_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_36_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_36_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_36_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_36_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_36_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_37_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_37_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_37_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_37_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_37_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_37_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_37_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_38_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_38_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_38_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_38_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_38_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_38_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_38_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_39_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_39_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_39_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_39_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_39_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_39_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_39_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_40_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_40_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_40_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_40_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_40_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_40_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_40_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_41_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_41_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_41_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_41_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_41_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_41_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_41_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_42_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_42_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_42_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_42_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_42_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_42_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_42_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_43_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_43_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_43_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_43_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_43_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_43_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_43_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_44_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_44_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_44_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_44_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_44_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_44_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_44_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_45_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_45_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_45_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_45_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_45_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_45_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_45_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_46_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_46_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_46_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_46_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_46_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_46_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_46_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_47_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_47_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_47_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_47_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_47_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_47_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_47_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_48_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_48_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_48_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_48_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_48_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_48_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_48_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_49_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_49_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_49_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_49_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_49_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_49_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_49_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_50_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_50_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_50_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_50_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_50_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_50_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_50_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_51_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_51_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_51_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_51_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_51_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_51_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_51_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_52_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_52_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_52_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_52_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_52_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_52_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_52_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_53_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_53_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_53_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_53_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_53_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_53_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_53_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_54_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_54_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_54_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_54_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_54_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_54_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_54_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_55_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_55_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_55_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_55_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_55_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_55_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_55_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_56_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_56_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_56_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_56_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_56_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_56_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_56_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_57_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_57_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_57_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_57_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_57_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_57_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_57_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_58_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_58_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_58_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_58_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_58_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_58_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_58_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_59_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_59_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_59_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_59_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_59_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_59_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_59_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_60_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_60_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_60_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_60_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_60_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_60_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_60_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_61_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_61_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_61_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_61_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_61_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_61_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_61_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_62_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_62_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_62_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_62_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_62_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_62_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_62_io_q0_next; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_63_io_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_63_io_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_63_io_q0; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_63_io_multiplicand; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_63_io_next_acc; // @[booth_multiplier.scala 23:33]
  wire [63:0] bs_63_io_next_Q; // @[booth_multiplier.scala 23:33]
  wire  bs_63_io_q0_next; // @[booth_multiplier.scala 23:33]
  booth_substep bs_0 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_0_io_acc),
    .io_Q(bs_0_io_Q),
    .io_q0(bs_0_io_q0),
    .io_multiplicand(bs_0_io_multiplicand),
    .io_next_acc(bs_0_io_next_acc),
    .io_next_Q(bs_0_io_next_Q),
    .io_q0_next(bs_0_io_q0_next)
  );
  booth_substep bs_1 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_1_io_acc),
    .io_Q(bs_1_io_Q),
    .io_q0(bs_1_io_q0),
    .io_multiplicand(bs_1_io_multiplicand),
    .io_next_acc(bs_1_io_next_acc),
    .io_next_Q(bs_1_io_next_Q),
    .io_q0_next(bs_1_io_q0_next)
  );
  booth_substep bs_2 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_2_io_acc),
    .io_Q(bs_2_io_Q),
    .io_q0(bs_2_io_q0),
    .io_multiplicand(bs_2_io_multiplicand),
    .io_next_acc(bs_2_io_next_acc),
    .io_next_Q(bs_2_io_next_Q),
    .io_q0_next(bs_2_io_q0_next)
  );
  booth_substep bs_3 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_3_io_acc),
    .io_Q(bs_3_io_Q),
    .io_q0(bs_3_io_q0),
    .io_multiplicand(bs_3_io_multiplicand),
    .io_next_acc(bs_3_io_next_acc),
    .io_next_Q(bs_3_io_next_Q),
    .io_q0_next(bs_3_io_q0_next)
  );
  booth_substep bs_4 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_4_io_acc),
    .io_Q(bs_4_io_Q),
    .io_q0(bs_4_io_q0),
    .io_multiplicand(bs_4_io_multiplicand),
    .io_next_acc(bs_4_io_next_acc),
    .io_next_Q(bs_4_io_next_Q),
    .io_q0_next(bs_4_io_q0_next)
  );
  booth_substep bs_5 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_5_io_acc),
    .io_Q(bs_5_io_Q),
    .io_q0(bs_5_io_q0),
    .io_multiplicand(bs_5_io_multiplicand),
    .io_next_acc(bs_5_io_next_acc),
    .io_next_Q(bs_5_io_next_Q),
    .io_q0_next(bs_5_io_q0_next)
  );
  booth_substep bs_6 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_6_io_acc),
    .io_Q(bs_6_io_Q),
    .io_q0(bs_6_io_q0),
    .io_multiplicand(bs_6_io_multiplicand),
    .io_next_acc(bs_6_io_next_acc),
    .io_next_Q(bs_6_io_next_Q),
    .io_q0_next(bs_6_io_q0_next)
  );
  booth_substep bs_7 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_7_io_acc),
    .io_Q(bs_7_io_Q),
    .io_q0(bs_7_io_q0),
    .io_multiplicand(bs_7_io_multiplicand),
    .io_next_acc(bs_7_io_next_acc),
    .io_next_Q(bs_7_io_next_Q),
    .io_q0_next(bs_7_io_q0_next)
  );
  booth_substep bs_8 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_8_io_acc),
    .io_Q(bs_8_io_Q),
    .io_q0(bs_8_io_q0),
    .io_multiplicand(bs_8_io_multiplicand),
    .io_next_acc(bs_8_io_next_acc),
    .io_next_Q(bs_8_io_next_Q),
    .io_q0_next(bs_8_io_q0_next)
  );
  booth_substep bs_9 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_9_io_acc),
    .io_Q(bs_9_io_Q),
    .io_q0(bs_9_io_q0),
    .io_multiplicand(bs_9_io_multiplicand),
    .io_next_acc(bs_9_io_next_acc),
    .io_next_Q(bs_9_io_next_Q),
    .io_q0_next(bs_9_io_q0_next)
  );
  booth_substep bs_10 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_10_io_acc),
    .io_Q(bs_10_io_Q),
    .io_q0(bs_10_io_q0),
    .io_multiplicand(bs_10_io_multiplicand),
    .io_next_acc(bs_10_io_next_acc),
    .io_next_Q(bs_10_io_next_Q),
    .io_q0_next(bs_10_io_q0_next)
  );
  booth_substep bs_11 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_11_io_acc),
    .io_Q(bs_11_io_Q),
    .io_q0(bs_11_io_q0),
    .io_multiplicand(bs_11_io_multiplicand),
    .io_next_acc(bs_11_io_next_acc),
    .io_next_Q(bs_11_io_next_Q),
    .io_q0_next(bs_11_io_q0_next)
  );
  booth_substep bs_12 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_12_io_acc),
    .io_Q(bs_12_io_Q),
    .io_q0(bs_12_io_q0),
    .io_multiplicand(bs_12_io_multiplicand),
    .io_next_acc(bs_12_io_next_acc),
    .io_next_Q(bs_12_io_next_Q),
    .io_q0_next(bs_12_io_q0_next)
  );
  booth_substep bs_13 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_13_io_acc),
    .io_Q(bs_13_io_Q),
    .io_q0(bs_13_io_q0),
    .io_multiplicand(bs_13_io_multiplicand),
    .io_next_acc(bs_13_io_next_acc),
    .io_next_Q(bs_13_io_next_Q),
    .io_q0_next(bs_13_io_q0_next)
  );
  booth_substep bs_14 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_14_io_acc),
    .io_Q(bs_14_io_Q),
    .io_q0(bs_14_io_q0),
    .io_multiplicand(bs_14_io_multiplicand),
    .io_next_acc(bs_14_io_next_acc),
    .io_next_Q(bs_14_io_next_Q),
    .io_q0_next(bs_14_io_q0_next)
  );
  booth_substep bs_15 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_15_io_acc),
    .io_Q(bs_15_io_Q),
    .io_q0(bs_15_io_q0),
    .io_multiplicand(bs_15_io_multiplicand),
    .io_next_acc(bs_15_io_next_acc),
    .io_next_Q(bs_15_io_next_Q),
    .io_q0_next(bs_15_io_q0_next)
  );
  booth_substep bs_16 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_16_io_acc),
    .io_Q(bs_16_io_Q),
    .io_q0(bs_16_io_q0),
    .io_multiplicand(bs_16_io_multiplicand),
    .io_next_acc(bs_16_io_next_acc),
    .io_next_Q(bs_16_io_next_Q),
    .io_q0_next(bs_16_io_q0_next)
  );
  booth_substep bs_17 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_17_io_acc),
    .io_Q(bs_17_io_Q),
    .io_q0(bs_17_io_q0),
    .io_multiplicand(bs_17_io_multiplicand),
    .io_next_acc(bs_17_io_next_acc),
    .io_next_Q(bs_17_io_next_Q),
    .io_q0_next(bs_17_io_q0_next)
  );
  booth_substep bs_18 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_18_io_acc),
    .io_Q(bs_18_io_Q),
    .io_q0(bs_18_io_q0),
    .io_multiplicand(bs_18_io_multiplicand),
    .io_next_acc(bs_18_io_next_acc),
    .io_next_Q(bs_18_io_next_Q),
    .io_q0_next(bs_18_io_q0_next)
  );
  booth_substep bs_19 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_19_io_acc),
    .io_Q(bs_19_io_Q),
    .io_q0(bs_19_io_q0),
    .io_multiplicand(bs_19_io_multiplicand),
    .io_next_acc(bs_19_io_next_acc),
    .io_next_Q(bs_19_io_next_Q),
    .io_q0_next(bs_19_io_q0_next)
  );
  booth_substep bs_20 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_20_io_acc),
    .io_Q(bs_20_io_Q),
    .io_q0(bs_20_io_q0),
    .io_multiplicand(bs_20_io_multiplicand),
    .io_next_acc(bs_20_io_next_acc),
    .io_next_Q(bs_20_io_next_Q),
    .io_q0_next(bs_20_io_q0_next)
  );
  booth_substep bs_21 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_21_io_acc),
    .io_Q(bs_21_io_Q),
    .io_q0(bs_21_io_q0),
    .io_multiplicand(bs_21_io_multiplicand),
    .io_next_acc(bs_21_io_next_acc),
    .io_next_Q(bs_21_io_next_Q),
    .io_q0_next(bs_21_io_q0_next)
  );
  booth_substep bs_22 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_22_io_acc),
    .io_Q(bs_22_io_Q),
    .io_q0(bs_22_io_q0),
    .io_multiplicand(bs_22_io_multiplicand),
    .io_next_acc(bs_22_io_next_acc),
    .io_next_Q(bs_22_io_next_Q),
    .io_q0_next(bs_22_io_q0_next)
  );
  booth_substep bs_23 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_23_io_acc),
    .io_Q(bs_23_io_Q),
    .io_q0(bs_23_io_q0),
    .io_multiplicand(bs_23_io_multiplicand),
    .io_next_acc(bs_23_io_next_acc),
    .io_next_Q(bs_23_io_next_Q),
    .io_q0_next(bs_23_io_q0_next)
  );
  booth_substep bs_24 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_24_io_acc),
    .io_Q(bs_24_io_Q),
    .io_q0(bs_24_io_q0),
    .io_multiplicand(bs_24_io_multiplicand),
    .io_next_acc(bs_24_io_next_acc),
    .io_next_Q(bs_24_io_next_Q),
    .io_q0_next(bs_24_io_q0_next)
  );
  booth_substep bs_25 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_25_io_acc),
    .io_Q(bs_25_io_Q),
    .io_q0(bs_25_io_q0),
    .io_multiplicand(bs_25_io_multiplicand),
    .io_next_acc(bs_25_io_next_acc),
    .io_next_Q(bs_25_io_next_Q),
    .io_q0_next(bs_25_io_q0_next)
  );
  booth_substep bs_26 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_26_io_acc),
    .io_Q(bs_26_io_Q),
    .io_q0(bs_26_io_q0),
    .io_multiplicand(bs_26_io_multiplicand),
    .io_next_acc(bs_26_io_next_acc),
    .io_next_Q(bs_26_io_next_Q),
    .io_q0_next(bs_26_io_q0_next)
  );
  booth_substep bs_27 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_27_io_acc),
    .io_Q(bs_27_io_Q),
    .io_q0(bs_27_io_q0),
    .io_multiplicand(bs_27_io_multiplicand),
    .io_next_acc(bs_27_io_next_acc),
    .io_next_Q(bs_27_io_next_Q),
    .io_q0_next(bs_27_io_q0_next)
  );
  booth_substep bs_28 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_28_io_acc),
    .io_Q(bs_28_io_Q),
    .io_q0(bs_28_io_q0),
    .io_multiplicand(bs_28_io_multiplicand),
    .io_next_acc(bs_28_io_next_acc),
    .io_next_Q(bs_28_io_next_Q),
    .io_q0_next(bs_28_io_q0_next)
  );
  booth_substep bs_29 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_29_io_acc),
    .io_Q(bs_29_io_Q),
    .io_q0(bs_29_io_q0),
    .io_multiplicand(bs_29_io_multiplicand),
    .io_next_acc(bs_29_io_next_acc),
    .io_next_Q(bs_29_io_next_Q),
    .io_q0_next(bs_29_io_q0_next)
  );
  booth_substep bs_30 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_30_io_acc),
    .io_Q(bs_30_io_Q),
    .io_q0(bs_30_io_q0),
    .io_multiplicand(bs_30_io_multiplicand),
    .io_next_acc(bs_30_io_next_acc),
    .io_next_Q(bs_30_io_next_Q),
    .io_q0_next(bs_30_io_q0_next)
  );
  booth_substep bs_31 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_31_io_acc),
    .io_Q(bs_31_io_Q),
    .io_q0(bs_31_io_q0),
    .io_multiplicand(bs_31_io_multiplicand),
    .io_next_acc(bs_31_io_next_acc),
    .io_next_Q(bs_31_io_next_Q),
    .io_q0_next(bs_31_io_q0_next)
  );
  booth_substep bs_32 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_32_io_acc),
    .io_Q(bs_32_io_Q),
    .io_q0(bs_32_io_q0),
    .io_multiplicand(bs_32_io_multiplicand),
    .io_next_acc(bs_32_io_next_acc),
    .io_next_Q(bs_32_io_next_Q),
    .io_q0_next(bs_32_io_q0_next)
  );
  booth_substep bs_33 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_33_io_acc),
    .io_Q(bs_33_io_Q),
    .io_q0(bs_33_io_q0),
    .io_multiplicand(bs_33_io_multiplicand),
    .io_next_acc(bs_33_io_next_acc),
    .io_next_Q(bs_33_io_next_Q),
    .io_q0_next(bs_33_io_q0_next)
  );
  booth_substep bs_34 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_34_io_acc),
    .io_Q(bs_34_io_Q),
    .io_q0(bs_34_io_q0),
    .io_multiplicand(bs_34_io_multiplicand),
    .io_next_acc(bs_34_io_next_acc),
    .io_next_Q(bs_34_io_next_Q),
    .io_q0_next(bs_34_io_q0_next)
  );
  booth_substep bs_35 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_35_io_acc),
    .io_Q(bs_35_io_Q),
    .io_q0(bs_35_io_q0),
    .io_multiplicand(bs_35_io_multiplicand),
    .io_next_acc(bs_35_io_next_acc),
    .io_next_Q(bs_35_io_next_Q),
    .io_q0_next(bs_35_io_q0_next)
  );
  booth_substep bs_36 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_36_io_acc),
    .io_Q(bs_36_io_Q),
    .io_q0(bs_36_io_q0),
    .io_multiplicand(bs_36_io_multiplicand),
    .io_next_acc(bs_36_io_next_acc),
    .io_next_Q(bs_36_io_next_Q),
    .io_q0_next(bs_36_io_q0_next)
  );
  booth_substep bs_37 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_37_io_acc),
    .io_Q(bs_37_io_Q),
    .io_q0(bs_37_io_q0),
    .io_multiplicand(bs_37_io_multiplicand),
    .io_next_acc(bs_37_io_next_acc),
    .io_next_Q(bs_37_io_next_Q),
    .io_q0_next(bs_37_io_q0_next)
  );
  booth_substep bs_38 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_38_io_acc),
    .io_Q(bs_38_io_Q),
    .io_q0(bs_38_io_q0),
    .io_multiplicand(bs_38_io_multiplicand),
    .io_next_acc(bs_38_io_next_acc),
    .io_next_Q(bs_38_io_next_Q),
    .io_q0_next(bs_38_io_q0_next)
  );
  booth_substep bs_39 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_39_io_acc),
    .io_Q(bs_39_io_Q),
    .io_q0(bs_39_io_q0),
    .io_multiplicand(bs_39_io_multiplicand),
    .io_next_acc(bs_39_io_next_acc),
    .io_next_Q(bs_39_io_next_Q),
    .io_q0_next(bs_39_io_q0_next)
  );
  booth_substep bs_40 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_40_io_acc),
    .io_Q(bs_40_io_Q),
    .io_q0(bs_40_io_q0),
    .io_multiplicand(bs_40_io_multiplicand),
    .io_next_acc(bs_40_io_next_acc),
    .io_next_Q(bs_40_io_next_Q),
    .io_q0_next(bs_40_io_q0_next)
  );
  booth_substep bs_41 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_41_io_acc),
    .io_Q(bs_41_io_Q),
    .io_q0(bs_41_io_q0),
    .io_multiplicand(bs_41_io_multiplicand),
    .io_next_acc(bs_41_io_next_acc),
    .io_next_Q(bs_41_io_next_Q),
    .io_q0_next(bs_41_io_q0_next)
  );
  booth_substep bs_42 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_42_io_acc),
    .io_Q(bs_42_io_Q),
    .io_q0(bs_42_io_q0),
    .io_multiplicand(bs_42_io_multiplicand),
    .io_next_acc(bs_42_io_next_acc),
    .io_next_Q(bs_42_io_next_Q),
    .io_q0_next(bs_42_io_q0_next)
  );
  booth_substep bs_43 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_43_io_acc),
    .io_Q(bs_43_io_Q),
    .io_q0(bs_43_io_q0),
    .io_multiplicand(bs_43_io_multiplicand),
    .io_next_acc(bs_43_io_next_acc),
    .io_next_Q(bs_43_io_next_Q),
    .io_q0_next(bs_43_io_q0_next)
  );
  booth_substep bs_44 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_44_io_acc),
    .io_Q(bs_44_io_Q),
    .io_q0(bs_44_io_q0),
    .io_multiplicand(bs_44_io_multiplicand),
    .io_next_acc(bs_44_io_next_acc),
    .io_next_Q(bs_44_io_next_Q),
    .io_q0_next(bs_44_io_q0_next)
  );
  booth_substep bs_45 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_45_io_acc),
    .io_Q(bs_45_io_Q),
    .io_q0(bs_45_io_q0),
    .io_multiplicand(bs_45_io_multiplicand),
    .io_next_acc(bs_45_io_next_acc),
    .io_next_Q(bs_45_io_next_Q),
    .io_q0_next(bs_45_io_q0_next)
  );
  booth_substep bs_46 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_46_io_acc),
    .io_Q(bs_46_io_Q),
    .io_q0(bs_46_io_q0),
    .io_multiplicand(bs_46_io_multiplicand),
    .io_next_acc(bs_46_io_next_acc),
    .io_next_Q(bs_46_io_next_Q),
    .io_q0_next(bs_46_io_q0_next)
  );
  booth_substep bs_47 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_47_io_acc),
    .io_Q(bs_47_io_Q),
    .io_q0(bs_47_io_q0),
    .io_multiplicand(bs_47_io_multiplicand),
    .io_next_acc(bs_47_io_next_acc),
    .io_next_Q(bs_47_io_next_Q),
    .io_q0_next(bs_47_io_q0_next)
  );
  booth_substep bs_48 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_48_io_acc),
    .io_Q(bs_48_io_Q),
    .io_q0(bs_48_io_q0),
    .io_multiplicand(bs_48_io_multiplicand),
    .io_next_acc(bs_48_io_next_acc),
    .io_next_Q(bs_48_io_next_Q),
    .io_q0_next(bs_48_io_q0_next)
  );
  booth_substep bs_49 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_49_io_acc),
    .io_Q(bs_49_io_Q),
    .io_q0(bs_49_io_q0),
    .io_multiplicand(bs_49_io_multiplicand),
    .io_next_acc(bs_49_io_next_acc),
    .io_next_Q(bs_49_io_next_Q),
    .io_q0_next(bs_49_io_q0_next)
  );
  booth_substep bs_50 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_50_io_acc),
    .io_Q(bs_50_io_Q),
    .io_q0(bs_50_io_q0),
    .io_multiplicand(bs_50_io_multiplicand),
    .io_next_acc(bs_50_io_next_acc),
    .io_next_Q(bs_50_io_next_Q),
    .io_q0_next(bs_50_io_q0_next)
  );
  booth_substep bs_51 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_51_io_acc),
    .io_Q(bs_51_io_Q),
    .io_q0(bs_51_io_q0),
    .io_multiplicand(bs_51_io_multiplicand),
    .io_next_acc(bs_51_io_next_acc),
    .io_next_Q(bs_51_io_next_Q),
    .io_q0_next(bs_51_io_q0_next)
  );
  booth_substep bs_52 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_52_io_acc),
    .io_Q(bs_52_io_Q),
    .io_q0(bs_52_io_q0),
    .io_multiplicand(bs_52_io_multiplicand),
    .io_next_acc(bs_52_io_next_acc),
    .io_next_Q(bs_52_io_next_Q),
    .io_q0_next(bs_52_io_q0_next)
  );
  booth_substep bs_53 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_53_io_acc),
    .io_Q(bs_53_io_Q),
    .io_q0(bs_53_io_q0),
    .io_multiplicand(bs_53_io_multiplicand),
    .io_next_acc(bs_53_io_next_acc),
    .io_next_Q(bs_53_io_next_Q),
    .io_q0_next(bs_53_io_q0_next)
  );
  booth_substep bs_54 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_54_io_acc),
    .io_Q(bs_54_io_Q),
    .io_q0(bs_54_io_q0),
    .io_multiplicand(bs_54_io_multiplicand),
    .io_next_acc(bs_54_io_next_acc),
    .io_next_Q(bs_54_io_next_Q),
    .io_q0_next(bs_54_io_q0_next)
  );
  booth_substep bs_55 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_55_io_acc),
    .io_Q(bs_55_io_Q),
    .io_q0(bs_55_io_q0),
    .io_multiplicand(bs_55_io_multiplicand),
    .io_next_acc(bs_55_io_next_acc),
    .io_next_Q(bs_55_io_next_Q),
    .io_q0_next(bs_55_io_q0_next)
  );
  booth_substep bs_56 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_56_io_acc),
    .io_Q(bs_56_io_Q),
    .io_q0(bs_56_io_q0),
    .io_multiplicand(bs_56_io_multiplicand),
    .io_next_acc(bs_56_io_next_acc),
    .io_next_Q(bs_56_io_next_Q),
    .io_q0_next(bs_56_io_q0_next)
  );
  booth_substep bs_57 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_57_io_acc),
    .io_Q(bs_57_io_Q),
    .io_q0(bs_57_io_q0),
    .io_multiplicand(bs_57_io_multiplicand),
    .io_next_acc(bs_57_io_next_acc),
    .io_next_Q(bs_57_io_next_Q),
    .io_q0_next(bs_57_io_q0_next)
  );
  booth_substep bs_58 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_58_io_acc),
    .io_Q(bs_58_io_Q),
    .io_q0(bs_58_io_q0),
    .io_multiplicand(bs_58_io_multiplicand),
    .io_next_acc(bs_58_io_next_acc),
    .io_next_Q(bs_58_io_next_Q),
    .io_q0_next(bs_58_io_q0_next)
  );
  booth_substep bs_59 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_59_io_acc),
    .io_Q(bs_59_io_Q),
    .io_q0(bs_59_io_q0),
    .io_multiplicand(bs_59_io_multiplicand),
    .io_next_acc(bs_59_io_next_acc),
    .io_next_Q(bs_59_io_next_Q),
    .io_q0_next(bs_59_io_q0_next)
  );
  booth_substep bs_60 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_60_io_acc),
    .io_Q(bs_60_io_Q),
    .io_q0(bs_60_io_q0),
    .io_multiplicand(bs_60_io_multiplicand),
    .io_next_acc(bs_60_io_next_acc),
    .io_next_Q(bs_60_io_next_Q),
    .io_q0_next(bs_60_io_q0_next)
  );
  booth_substep bs_61 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_61_io_acc),
    .io_Q(bs_61_io_Q),
    .io_q0(bs_61_io_q0),
    .io_multiplicand(bs_61_io_multiplicand),
    .io_next_acc(bs_61_io_next_acc),
    .io_next_Q(bs_61_io_next_Q),
    .io_q0_next(bs_61_io_q0_next)
  );
  booth_substep bs_62 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_62_io_acc),
    .io_Q(bs_62_io_Q),
    .io_q0(bs_62_io_q0),
    .io_multiplicand(bs_62_io_multiplicand),
    .io_next_acc(bs_62_io_next_acc),
    .io_next_Q(bs_62_io_next_Q),
    .io_q0_next(bs_62_io_q0_next)
  );
  booth_substep bs_63 ( // @[booth_multiplier.scala 23:33]
    .io_acc(bs_63_io_acc),
    .io_Q(bs_63_io_Q),
    .io_q0(bs_63_io_q0),
    .io_multiplicand(bs_63_io_multiplicand),
    .io_next_acc(bs_63_io_next_acc),
    .io_next_Q(bs_63_io_next_Q),
    .io_q0_next(bs_63_io_q0_next)
  );
  assign io_product = {bs_63_io_next_acc,bs_63_io_next_Q}; // @[booth_multiplier.scala 43:56]
  assign bs_0_io_acc = 64'sh0; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 20:12]
  assign bs_0_io_Q = io_multiplier; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 21:10]
  assign bs_0_io_q0 = 1'h0; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 19:11]
  assign bs_0_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_1_io_acc = bs_0_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_1_io_Q = bs_0_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_1_io_q0 = bs_0_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_1_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_2_io_acc = bs_1_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_2_io_Q = bs_1_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_2_io_q0 = bs_1_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_2_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_3_io_acc = bs_2_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_3_io_Q = bs_2_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_3_io_q0 = bs_2_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_3_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_4_io_acc = bs_3_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_4_io_Q = bs_3_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_4_io_q0 = bs_3_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_4_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_5_io_acc = bs_4_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_5_io_Q = bs_4_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_5_io_q0 = bs_4_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_5_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_6_io_acc = bs_5_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_6_io_Q = bs_5_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_6_io_q0 = bs_5_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_6_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_7_io_acc = bs_6_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_7_io_Q = bs_6_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_7_io_q0 = bs_6_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_7_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_8_io_acc = bs_7_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_8_io_Q = bs_7_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_8_io_q0 = bs_7_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_8_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_9_io_acc = bs_8_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_9_io_Q = bs_8_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_9_io_q0 = bs_8_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_9_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_10_io_acc = bs_9_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_10_io_Q = bs_9_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_10_io_q0 = bs_9_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_10_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_11_io_acc = bs_10_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_11_io_Q = bs_10_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_11_io_q0 = bs_10_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_11_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_12_io_acc = bs_11_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_12_io_Q = bs_11_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_12_io_q0 = bs_11_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_12_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_13_io_acc = bs_12_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_13_io_Q = bs_12_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_13_io_q0 = bs_12_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_13_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_14_io_acc = bs_13_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_14_io_Q = bs_13_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_14_io_q0 = bs_13_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_14_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_15_io_acc = bs_14_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_15_io_Q = bs_14_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_15_io_q0 = bs_14_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_15_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_16_io_acc = bs_15_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_16_io_Q = bs_15_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_16_io_q0 = bs_15_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_16_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_17_io_acc = bs_16_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_17_io_Q = bs_16_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_17_io_q0 = bs_16_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_17_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_18_io_acc = bs_17_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_18_io_Q = bs_17_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_18_io_q0 = bs_17_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_18_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_19_io_acc = bs_18_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_19_io_Q = bs_18_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_19_io_q0 = bs_18_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_19_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_20_io_acc = bs_19_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_20_io_Q = bs_19_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_20_io_q0 = bs_19_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_20_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_21_io_acc = bs_20_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_21_io_Q = bs_20_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_21_io_q0 = bs_20_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_21_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_22_io_acc = bs_21_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_22_io_Q = bs_21_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_22_io_q0 = bs_21_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_22_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_23_io_acc = bs_22_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_23_io_Q = bs_22_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_23_io_q0 = bs_22_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_23_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_24_io_acc = bs_23_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_24_io_Q = bs_23_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_24_io_q0 = bs_23_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_24_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_25_io_acc = bs_24_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_25_io_Q = bs_24_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_25_io_q0 = bs_24_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_25_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_26_io_acc = bs_25_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_26_io_Q = bs_25_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_26_io_q0 = bs_25_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_26_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_27_io_acc = bs_26_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_27_io_Q = bs_26_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_27_io_q0 = bs_26_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_27_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_28_io_acc = bs_27_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_28_io_Q = bs_27_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_28_io_q0 = bs_27_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_28_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_29_io_acc = bs_28_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_29_io_Q = bs_28_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_29_io_q0 = bs_28_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_29_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_30_io_acc = bs_29_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_30_io_Q = bs_29_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_30_io_q0 = bs_29_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_30_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_31_io_acc = bs_30_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_31_io_Q = bs_30_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_31_io_q0 = bs_30_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_31_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_32_io_acc = bs_31_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_32_io_Q = bs_31_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_32_io_q0 = bs_31_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_32_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_33_io_acc = bs_32_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_33_io_Q = bs_32_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_33_io_q0 = bs_32_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_33_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_34_io_acc = bs_33_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_34_io_Q = bs_33_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_34_io_q0 = bs_33_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_34_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_35_io_acc = bs_34_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_35_io_Q = bs_34_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_35_io_q0 = bs_34_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_35_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_36_io_acc = bs_35_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_36_io_Q = bs_35_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_36_io_q0 = bs_35_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_36_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_37_io_acc = bs_36_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_37_io_Q = bs_36_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_37_io_q0 = bs_36_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_37_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_38_io_acc = bs_37_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_38_io_Q = bs_37_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_38_io_q0 = bs_37_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_38_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_39_io_acc = bs_38_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_39_io_Q = bs_38_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_39_io_q0 = bs_38_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_39_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_40_io_acc = bs_39_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_40_io_Q = bs_39_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_40_io_q0 = bs_39_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_40_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_41_io_acc = bs_40_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_41_io_Q = bs_40_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_41_io_q0 = bs_40_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_41_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_42_io_acc = bs_41_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_42_io_Q = bs_41_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_42_io_q0 = bs_41_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_42_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_43_io_acc = bs_42_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_43_io_Q = bs_42_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_43_io_q0 = bs_42_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_43_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_44_io_acc = bs_43_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_44_io_Q = bs_43_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_44_io_q0 = bs_43_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_44_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_45_io_acc = bs_44_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_45_io_Q = bs_44_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_45_io_q0 = bs_44_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_45_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_46_io_acc = bs_45_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_46_io_Q = bs_45_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_46_io_q0 = bs_45_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_46_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_47_io_acc = bs_46_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_47_io_Q = bs_46_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_47_io_q0 = bs_46_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_47_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_48_io_acc = bs_47_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_48_io_Q = bs_47_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_48_io_q0 = bs_47_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_48_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_49_io_acc = bs_48_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_49_io_Q = bs_48_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_49_io_q0 = bs_48_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_49_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_50_io_acc = bs_49_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_50_io_Q = bs_49_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_50_io_q0 = bs_49_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_50_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_51_io_acc = bs_50_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_51_io_Q = bs_50_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_51_io_q0 = bs_50_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_51_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_52_io_acc = bs_51_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_52_io_Q = bs_51_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_52_io_q0 = bs_51_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_52_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_53_io_acc = bs_52_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_53_io_Q = bs_52_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_53_io_q0 = bs_52_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_53_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_54_io_acc = bs_53_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_54_io_Q = bs_53_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_54_io_q0 = bs_53_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_54_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_55_io_acc = bs_54_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_55_io_Q = bs_54_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_55_io_q0 = bs_54_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_55_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_56_io_acc = bs_55_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_56_io_Q = bs_55_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_56_io_q0 = bs_55_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_56_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_57_io_acc = bs_56_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_57_io_Q = bs_56_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_57_io_q0 = bs_56_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_57_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_58_io_acc = bs_57_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_58_io_Q = bs_57_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_58_io_q0 = bs_57_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_58_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_59_io_acc = bs_58_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_59_io_Q = bs_58_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_59_io_q0 = bs_58_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_59_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_60_io_acc = bs_59_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_60_io_Q = bs_59_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_60_io_q0 = bs_59_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_60_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_61_io_acc = bs_60_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_61_io_Q = bs_60_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_61_io_q0 = bs_60_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_61_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_62_io_acc = bs_61_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_62_io_Q = bs_61_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_62_io_q0 = bs_61_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_62_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 29:31]
  assign bs_63_io_acc = bs_62_io_next_acc; // @[booth_multiplier.scala 12:19 booth_multiplier.scala 30:18]
  assign bs_63_io_Q = bs_62_io_next_Q; // @[booth_multiplier.scala 11:17 booth_multiplier.scala 31:16]
  assign bs_63_io_q0 = bs_62_io_q0_next; // @[booth_multiplier.scala 13:18 booth_multiplier.scala 32:17]
  assign bs_63_io_multiplicand = io_multiplicand; // @[booth_multiplier.scala 38:28]
endmodule
