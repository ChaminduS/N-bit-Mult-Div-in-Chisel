module fullAdder(
  input   io_i0,
  input   io_i1,
  input   io_cin,
  output  io_sum,
  output  io_cout
);
  assign io_sum = io_i0 ^ io_i1 ^ io_cin; // @[addsub_64.scala 14:29]
  assign io_cout = io_i0 & io_i1 | io_i1 & io_cin | io_cin & io_i0; // @[addsub_64.scala 15:51]
endmodule
module addsub_64(
  input         clock,
  input         reset,
  input         io_cin,
  input  [63:0] io_onesComp_ip,
  input  [63:0] io_i0,
  output [63:0] io_sum
);
  wire  fa_0_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_0_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_0_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_0_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_0_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_1_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_1_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_1_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_1_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_1_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_2_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_2_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_2_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_2_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_2_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_3_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_3_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_3_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_3_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_3_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_4_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_4_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_4_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_4_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_4_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_5_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_5_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_5_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_5_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_5_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_6_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_6_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_6_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_6_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_6_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_7_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_7_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_7_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_7_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_7_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_8_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_8_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_8_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_8_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_8_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_9_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_9_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_9_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_9_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_9_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_10_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_10_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_10_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_10_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_10_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_11_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_11_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_11_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_11_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_11_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_12_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_12_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_12_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_12_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_12_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_13_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_13_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_13_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_13_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_13_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_14_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_14_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_14_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_14_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_14_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_15_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_15_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_15_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_15_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_15_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_16_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_16_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_16_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_16_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_16_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_17_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_17_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_17_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_17_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_17_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_18_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_18_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_18_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_18_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_18_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_19_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_19_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_19_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_19_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_19_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_20_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_20_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_20_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_20_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_20_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_21_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_21_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_21_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_21_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_21_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_22_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_22_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_22_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_22_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_22_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_23_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_23_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_23_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_23_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_23_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_24_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_24_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_24_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_24_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_24_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_25_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_25_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_25_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_25_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_25_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_26_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_26_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_26_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_26_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_26_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_27_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_27_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_27_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_27_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_27_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_28_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_28_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_28_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_28_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_28_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_29_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_29_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_29_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_29_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_29_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_30_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_30_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_30_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_30_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_30_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_31_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_31_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_31_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_31_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_31_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_32_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_32_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_32_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_32_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_32_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_33_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_33_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_33_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_33_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_33_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_34_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_34_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_34_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_34_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_34_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_35_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_35_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_35_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_35_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_35_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_36_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_36_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_36_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_36_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_36_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_37_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_37_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_37_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_37_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_37_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_38_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_38_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_38_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_38_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_38_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_39_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_39_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_39_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_39_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_39_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_40_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_40_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_40_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_40_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_40_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_41_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_41_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_41_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_41_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_41_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_42_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_42_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_42_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_42_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_42_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_43_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_43_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_43_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_43_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_43_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_44_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_44_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_44_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_44_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_44_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_45_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_45_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_45_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_45_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_45_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_46_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_46_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_46_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_46_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_46_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_47_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_47_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_47_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_47_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_47_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_48_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_48_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_48_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_48_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_48_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_49_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_49_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_49_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_49_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_49_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_50_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_50_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_50_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_50_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_50_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_51_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_51_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_51_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_51_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_51_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_52_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_52_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_52_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_52_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_52_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_53_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_53_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_53_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_53_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_53_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_54_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_54_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_54_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_54_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_54_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_55_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_55_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_55_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_55_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_55_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_56_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_56_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_56_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_56_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_56_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_57_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_57_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_57_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_57_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_57_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_58_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_58_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_58_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_58_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_58_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_59_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_59_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_59_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_59_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_59_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_60_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_60_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_60_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_60_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_60_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_61_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_61_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_61_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_61_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_61_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_62_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_62_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_62_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_62_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_62_io_cout; // @[addsub_64.scala 27:33]
  wire  fa_63_io_i0; // @[addsub_64.scala 27:33]
  wire  fa_63_io_i1; // @[addsub_64.scala 27:33]
  wire  fa_63_io_cin; // @[addsub_64.scala 27:33]
  wire  fa_63_io_sum; // @[addsub_64.scala 27:33]
  wire  fa_63_io_cout; // @[addsub_64.scala 27:33]
  wire [7:0] lo_lo_lo = {fa_7_io_sum,fa_6_io_sum,fa_5_io_sum,fa_4_io_sum,fa_3_io_sum,fa_2_io_sum,fa_1_io_sum,fa_0_io_sum
    }; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {fa_15_io_sum,fa_14_io_sum,fa_13_io_sum,fa_12_io_sum,fa_11_io_sum,fa_10_io_sum,fa_9_io_sum,
    fa_8_io_sum,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {fa_23_io_sum,fa_22_io_sum,fa_21_io_sum,fa_20_io_sum,fa_19_io_sum,fa_18_io_sum,fa_17_io_sum,
    fa_16_io_sum}; // @[Cat.scala 30:58]
  wire [31:0] lo = {fa_31_io_sum,fa_30_io_sum,fa_29_io_sum,fa_28_io_sum,fa_27_io_sum,fa_26_io_sum,fa_25_io_sum,
    fa_24_io_sum,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {fa_39_io_sum,fa_38_io_sum,fa_37_io_sum,fa_36_io_sum,fa_35_io_sum,fa_34_io_sum,fa_33_io_sum,
    fa_32_io_sum}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {fa_47_io_sum,fa_46_io_sum,fa_45_io_sum,fa_44_io_sum,fa_43_io_sum,fa_42_io_sum,fa_41_io_sum,
    fa_40_io_sum,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {fa_55_io_sum,fa_54_io_sum,fa_53_io_sum,fa_52_io_sum,fa_51_io_sum,fa_50_io_sum,fa_49_io_sum,
    fa_48_io_sum}; // @[Cat.scala 30:58]
  wire [31:0] hi = {fa_63_io_sum,fa_62_io_sum,fa_61_io_sum,fa_60_io_sum,fa_59_io_sum,fa_58_io_sum,fa_57_io_sum,
    fa_56_io_sum,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  fullAdder fa_0 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_0_io_i0),
    .io_i1(fa_0_io_i1),
    .io_cin(fa_0_io_cin),
    .io_sum(fa_0_io_sum),
    .io_cout(fa_0_io_cout)
  );
  fullAdder fa_1 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_1_io_i0),
    .io_i1(fa_1_io_i1),
    .io_cin(fa_1_io_cin),
    .io_sum(fa_1_io_sum),
    .io_cout(fa_1_io_cout)
  );
  fullAdder fa_2 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_2_io_i0),
    .io_i1(fa_2_io_i1),
    .io_cin(fa_2_io_cin),
    .io_sum(fa_2_io_sum),
    .io_cout(fa_2_io_cout)
  );
  fullAdder fa_3 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_3_io_i0),
    .io_i1(fa_3_io_i1),
    .io_cin(fa_3_io_cin),
    .io_sum(fa_3_io_sum),
    .io_cout(fa_3_io_cout)
  );
  fullAdder fa_4 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_4_io_i0),
    .io_i1(fa_4_io_i1),
    .io_cin(fa_4_io_cin),
    .io_sum(fa_4_io_sum),
    .io_cout(fa_4_io_cout)
  );
  fullAdder fa_5 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_5_io_i0),
    .io_i1(fa_5_io_i1),
    .io_cin(fa_5_io_cin),
    .io_sum(fa_5_io_sum),
    .io_cout(fa_5_io_cout)
  );
  fullAdder fa_6 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_6_io_i0),
    .io_i1(fa_6_io_i1),
    .io_cin(fa_6_io_cin),
    .io_sum(fa_6_io_sum),
    .io_cout(fa_6_io_cout)
  );
  fullAdder fa_7 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_7_io_i0),
    .io_i1(fa_7_io_i1),
    .io_cin(fa_7_io_cin),
    .io_sum(fa_7_io_sum),
    .io_cout(fa_7_io_cout)
  );
  fullAdder fa_8 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_8_io_i0),
    .io_i1(fa_8_io_i1),
    .io_cin(fa_8_io_cin),
    .io_sum(fa_8_io_sum),
    .io_cout(fa_8_io_cout)
  );
  fullAdder fa_9 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_9_io_i0),
    .io_i1(fa_9_io_i1),
    .io_cin(fa_9_io_cin),
    .io_sum(fa_9_io_sum),
    .io_cout(fa_9_io_cout)
  );
  fullAdder fa_10 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_10_io_i0),
    .io_i1(fa_10_io_i1),
    .io_cin(fa_10_io_cin),
    .io_sum(fa_10_io_sum),
    .io_cout(fa_10_io_cout)
  );
  fullAdder fa_11 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_11_io_i0),
    .io_i1(fa_11_io_i1),
    .io_cin(fa_11_io_cin),
    .io_sum(fa_11_io_sum),
    .io_cout(fa_11_io_cout)
  );
  fullAdder fa_12 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_12_io_i0),
    .io_i1(fa_12_io_i1),
    .io_cin(fa_12_io_cin),
    .io_sum(fa_12_io_sum),
    .io_cout(fa_12_io_cout)
  );
  fullAdder fa_13 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_13_io_i0),
    .io_i1(fa_13_io_i1),
    .io_cin(fa_13_io_cin),
    .io_sum(fa_13_io_sum),
    .io_cout(fa_13_io_cout)
  );
  fullAdder fa_14 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_14_io_i0),
    .io_i1(fa_14_io_i1),
    .io_cin(fa_14_io_cin),
    .io_sum(fa_14_io_sum),
    .io_cout(fa_14_io_cout)
  );
  fullAdder fa_15 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_15_io_i0),
    .io_i1(fa_15_io_i1),
    .io_cin(fa_15_io_cin),
    .io_sum(fa_15_io_sum),
    .io_cout(fa_15_io_cout)
  );
  fullAdder fa_16 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_16_io_i0),
    .io_i1(fa_16_io_i1),
    .io_cin(fa_16_io_cin),
    .io_sum(fa_16_io_sum),
    .io_cout(fa_16_io_cout)
  );
  fullAdder fa_17 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_17_io_i0),
    .io_i1(fa_17_io_i1),
    .io_cin(fa_17_io_cin),
    .io_sum(fa_17_io_sum),
    .io_cout(fa_17_io_cout)
  );
  fullAdder fa_18 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_18_io_i0),
    .io_i1(fa_18_io_i1),
    .io_cin(fa_18_io_cin),
    .io_sum(fa_18_io_sum),
    .io_cout(fa_18_io_cout)
  );
  fullAdder fa_19 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_19_io_i0),
    .io_i1(fa_19_io_i1),
    .io_cin(fa_19_io_cin),
    .io_sum(fa_19_io_sum),
    .io_cout(fa_19_io_cout)
  );
  fullAdder fa_20 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_20_io_i0),
    .io_i1(fa_20_io_i1),
    .io_cin(fa_20_io_cin),
    .io_sum(fa_20_io_sum),
    .io_cout(fa_20_io_cout)
  );
  fullAdder fa_21 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_21_io_i0),
    .io_i1(fa_21_io_i1),
    .io_cin(fa_21_io_cin),
    .io_sum(fa_21_io_sum),
    .io_cout(fa_21_io_cout)
  );
  fullAdder fa_22 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_22_io_i0),
    .io_i1(fa_22_io_i1),
    .io_cin(fa_22_io_cin),
    .io_sum(fa_22_io_sum),
    .io_cout(fa_22_io_cout)
  );
  fullAdder fa_23 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_23_io_i0),
    .io_i1(fa_23_io_i1),
    .io_cin(fa_23_io_cin),
    .io_sum(fa_23_io_sum),
    .io_cout(fa_23_io_cout)
  );
  fullAdder fa_24 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_24_io_i0),
    .io_i1(fa_24_io_i1),
    .io_cin(fa_24_io_cin),
    .io_sum(fa_24_io_sum),
    .io_cout(fa_24_io_cout)
  );
  fullAdder fa_25 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_25_io_i0),
    .io_i1(fa_25_io_i1),
    .io_cin(fa_25_io_cin),
    .io_sum(fa_25_io_sum),
    .io_cout(fa_25_io_cout)
  );
  fullAdder fa_26 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_26_io_i0),
    .io_i1(fa_26_io_i1),
    .io_cin(fa_26_io_cin),
    .io_sum(fa_26_io_sum),
    .io_cout(fa_26_io_cout)
  );
  fullAdder fa_27 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_27_io_i0),
    .io_i1(fa_27_io_i1),
    .io_cin(fa_27_io_cin),
    .io_sum(fa_27_io_sum),
    .io_cout(fa_27_io_cout)
  );
  fullAdder fa_28 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_28_io_i0),
    .io_i1(fa_28_io_i1),
    .io_cin(fa_28_io_cin),
    .io_sum(fa_28_io_sum),
    .io_cout(fa_28_io_cout)
  );
  fullAdder fa_29 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_29_io_i0),
    .io_i1(fa_29_io_i1),
    .io_cin(fa_29_io_cin),
    .io_sum(fa_29_io_sum),
    .io_cout(fa_29_io_cout)
  );
  fullAdder fa_30 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_30_io_i0),
    .io_i1(fa_30_io_i1),
    .io_cin(fa_30_io_cin),
    .io_sum(fa_30_io_sum),
    .io_cout(fa_30_io_cout)
  );
  fullAdder fa_31 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_31_io_i0),
    .io_i1(fa_31_io_i1),
    .io_cin(fa_31_io_cin),
    .io_sum(fa_31_io_sum),
    .io_cout(fa_31_io_cout)
  );
  fullAdder fa_32 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_32_io_i0),
    .io_i1(fa_32_io_i1),
    .io_cin(fa_32_io_cin),
    .io_sum(fa_32_io_sum),
    .io_cout(fa_32_io_cout)
  );
  fullAdder fa_33 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_33_io_i0),
    .io_i1(fa_33_io_i1),
    .io_cin(fa_33_io_cin),
    .io_sum(fa_33_io_sum),
    .io_cout(fa_33_io_cout)
  );
  fullAdder fa_34 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_34_io_i0),
    .io_i1(fa_34_io_i1),
    .io_cin(fa_34_io_cin),
    .io_sum(fa_34_io_sum),
    .io_cout(fa_34_io_cout)
  );
  fullAdder fa_35 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_35_io_i0),
    .io_i1(fa_35_io_i1),
    .io_cin(fa_35_io_cin),
    .io_sum(fa_35_io_sum),
    .io_cout(fa_35_io_cout)
  );
  fullAdder fa_36 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_36_io_i0),
    .io_i1(fa_36_io_i1),
    .io_cin(fa_36_io_cin),
    .io_sum(fa_36_io_sum),
    .io_cout(fa_36_io_cout)
  );
  fullAdder fa_37 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_37_io_i0),
    .io_i1(fa_37_io_i1),
    .io_cin(fa_37_io_cin),
    .io_sum(fa_37_io_sum),
    .io_cout(fa_37_io_cout)
  );
  fullAdder fa_38 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_38_io_i0),
    .io_i1(fa_38_io_i1),
    .io_cin(fa_38_io_cin),
    .io_sum(fa_38_io_sum),
    .io_cout(fa_38_io_cout)
  );
  fullAdder fa_39 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_39_io_i0),
    .io_i1(fa_39_io_i1),
    .io_cin(fa_39_io_cin),
    .io_sum(fa_39_io_sum),
    .io_cout(fa_39_io_cout)
  );
  fullAdder fa_40 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_40_io_i0),
    .io_i1(fa_40_io_i1),
    .io_cin(fa_40_io_cin),
    .io_sum(fa_40_io_sum),
    .io_cout(fa_40_io_cout)
  );
  fullAdder fa_41 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_41_io_i0),
    .io_i1(fa_41_io_i1),
    .io_cin(fa_41_io_cin),
    .io_sum(fa_41_io_sum),
    .io_cout(fa_41_io_cout)
  );
  fullAdder fa_42 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_42_io_i0),
    .io_i1(fa_42_io_i1),
    .io_cin(fa_42_io_cin),
    .io_sum(fa_42_io_sum),
    .io_cout(fa_42_io_cout)
  );
  fullAdder fa_43 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_43_io_i0),
    .io_i1(fa_43_io_i1),
    .io_cin(fa_43_io_cin),
    .io_sum(fa_43_io_sum),
    .io_cout(fa_43_io_cout)
  );
  fullAdder fa_44 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_44_io_i0),
    .io_i1(fa_44_io_i1),
    .io_cin(fa_44_io_cin),
    .io_sum(fa_44_io_sum),
    .io_cout(fa_44_io_cout)
  );
  fullAdder fa_45 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_45_io_i0),
    .io_i1(fa_45_io_i1),
    .io_cin(fa_45_io_cin),
    .io_sum(fa_45_io_sum),
    .io_cout(fa_45_io_cout)
  );
  fullAdder fa_46 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_46_io_i0),
    .io_i1(fa_46_io_i1),
    .io_cin(fa_46_io_cin),
    .io_sum(fa_46_io_sum),
    .io_cout(fa_46_io_cout)
  );
  fullAdder fa_47 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_47_io_i0),
    .io_i1(fa_47_io_i1),
    .io_cin(fa_47_io_cin),
    .io_sum(fa_47_io_sum),
    .io_cout(fa_47_io_cout)
  );
  fullAdder fa_48 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_48_io_i0),
    .io_i1(fa_48_io_i1),
    .io_cin(fa_48_io_cin),
    .io_sum(fa_48_io_sum),
    .io_cout(fa_48_io_cout)
  );
  fullAdder fa_49 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_49_io_i0),
    .io_i1(fa_49_io_i1),
    .io_cin(fa_49_io_cin),
    .io_sum(fa_49_io_sum),
    .io_cout(fa_49_io_cout)
  );
  fullAdder fa_50 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_50_io_i0),
    .io_i1(fa_50_io_i1),
    .io_cin(fa_50_io_cin),
    .io_sum(fa_50_io_sum),
    .io_cout(fa_50_io_cout)
  );
  fullAdder fa_51 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_51_io_i0),
    .io_i1(fa_51_io_i1),
    .io_cin(fa_51_io_cin),
    .io_sum(fa_51_io_sum),
    .io_cout(fa_51_io_cout)
  );
  fullAdder fa_52 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_52_io_i0),
    .io_i1(fa_52_io_i1),
    .io_cin(fa_52_io_cin),
    .io_sum(fa_52_io_sum),
    .io_cout(fa_52_io_cout)
  );
  fullAdder fa_53 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_53_io_i0),
    .io_i1(fa_53_io_i1),
    .io_cin(fa_53_io_cin),
    .io_sum(fa_53_io_sum),
    .io_cout(fa_53_io_cout)
  );
  fullAdder fa_54 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_54_io_i0),
    .io_i1(fa_54_io_i1),
    .io_cin(fa_54_io_cin),
    .io_sum(fa_54_io_sum),
    .io_cout(fa_54_io_cout)
  );
  fullAdder fa_55 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_55_io_i0),
    .io_i1(fa_55_io_i1),
    .io_cin(fa_55_io_cin),
    .io_sum(fa_55_io_sum),
    .io_cout(fa_55_io_cout)
  );
  fullAdder fa_56 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_56_io_i0),
    .io_i1(fa_56_io_i1),
    .io_cin(fa_56_io_cin),
    .io_sum(fa_56_io_sum),
    .io_cout(fa_56_io_cout)
  );
  fullAdder fa_57 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_57_io_i0),
    .io_i1(fa_57_io_i1),
    .io_cin(fa_57_io_cin),
    .io_sum(fa_57_io_sum),
    .io_cout(fa_57_io_cout)
  );
  fullAdder fa_58 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_58_io_i0),
    .io_i1(fa_58_io_i1),
    .io_cin(fa_58_io_cin),
    .io_sum(fa_58_io_sum),
    .io_cout(fa_58_io_cout)
  );
  fullAdder fa_59 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_59_io_i0),
    .io_i1(fa_59_io_i1),
    .io_cin(fa_59_io_cin),
    .io_sum(fa_59_io_sum),
    .io_cout(fa_59_io_cout)
  );
  fullAdder fa_60 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_60_io_i0),
    .io_i1(fa_60_io_i1),
    .io_cin(fa_60_io_cin),
    .io_sum(fa_60_io_sum),
    .io_cout(fa_60_io_cout)
  );
  fullAdder fa_61 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_61_io_i0),
    .io_i1(fa_61_io_i1),
    .io_cin(fa_61_io_cin),
    .io_sum(fa_61_io_sum),
    .io_cout(fa_61_io_cout)
  );
  fullAdder fa_62 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_62_io_i0),
    .io_i1(fa_62_io_i1),
    .io_cin(fa_62_io_cin),
    .io_sum(fa_62_io_sum),
    .io_cout(fa_62_io_cout)
  );
  fullAdder fa_63 ( // @[addsub_64.scala 27:33]
    .io_i0(fa_63_io_i0),
    .io_i1(fa_63_io_i1),
    .io_cin(fa_63_io_cin),
    .io_sum(fa_63_io_sum),
    .io_cout(fa_63_io_cout)
  );
  assign io_sum = {hi,lo}; // @[Cat.scala 30:58]
  assign fa_0_io_i0 = io_i0[0]; // @[addsub_64.scala 31:25]
  assign fa_0_io_i1 = io_onesComp_ip[0]; // @[addsub_64.scala 32:34]
  assign fa_0_io_cin = io_cin; // @[addsub_64.scala 33:18]
  assign fa_1_io_i0 = io_i0[1]; // @[addsub_64.scala 37:29]
  assign fa_1_io_i1 = io_onesComp_ip[1]; // @[addsub_64.scala 38:38]
  assign fa_1_io_cin = fa_0_io_cout; // @[addsub_64.scala 39:22]
  assign fa_2_io_i0 = io_i0[2]; // @[addsub_64.scala 37:29]
  assign fa_2_io_i1 = io_onesComp_ip[2]; // @[addsub_64.scala 38:38]
  assign fa_2_io_cin = fa_1_io_cout; // @[addsub_64.scala 39:22]
  assign fa_3_io_i0 = io_i0[3]; // @[addsub_64.scala 37:29]
  assign fa_3_io_i1 = io_onesComp_ip[3]; // @[addsub_64.scala 38:38]
  assign fa_3_io_cin = fa_2_io_cout; // @[addsub_64.scala 39:22]
  assign fa_4_io_i0 = io_i0[4]; // @[addsub_64.scala 37:29]
  assign fa_4_io_i1 = io_onesComp_ip[4]; // @[addsub_64.scala 38:38]
  assign fa_4_io_cin = fa_3_io_cout; // @[addsub_64.scala 39:22]
  assign fa_5_io_i0 = io_i0[5]; // @[addsub_64.scala 37:29]
  assign fa_5_io_i1 = io_onesComp_ip[5]; // @[addsub_64.scala 38:38]
  assign fa_5_io_cin = fa_4_io_cout; // @[addsub_64.scala 39:22]
  assign fa_6_io_i0 = io_i0[6]; // @[addsub_64.scala 37:29]
  assign fa_6_io_i1 = io_onesComp_ip[6]; // @[addsub_64.scala 38:38]
  assign fa_6_io_cin = fa_5_io_cout; // @[addsub_64.scala 39:22]
  assign fa_7_io_i0 = io_i0[7]; // @[addsub_64.scala 37:29]
  assign fa_7_io_i1 = io_onesComp_ip[7]; // @[addsub_64.scala 38:38]
  assign fa_7_io_cin = fa_6_io_cout; // @[addsub_64.scala 39:22]
  assign fa_8_io_i0 = io_i0[8]; // @[addsub_64.scala 37:29]
  assign fa_8_io_i1 = io_onesComp_ip[8]; // @[addsub_64.scala 38:38]
  assign fa_8_io_cin = fa_7_io_cout; // @[addsub_64.scala 39:22]
  assign fa_9_io_i0 = io_i0[9]; // @[addsub_64.scala 37:29]
  assign fa_9_io_i1 = io_onesComp_ip[9]; // @[addsub_64.scala 38:38]
  assign fa_9_io_cin = fa_8_io_cout; // @[addsub_64.scala 39:22]
  assign fa_10_io_i0 = io_i0[10]; // @[addsub_64.scala 37:29]
  assign fa_10_io_i1 = io_onesComp_ip[10]; // @[addsub_64.scala 38:38]
  assign fa_10_io_cin = fa_9_io_cout; // @[addsub_64.scala 39:22]
  assign fa_11_io_i0 = io_i0[11]; // @[addsub_64.scala 37:29]
  assign fa_11_io_i1 = io_onesComp_ip[11]; // @[addsub_64.scala 38:38]
  assign fa_11_io_cin = fa_10_io_cout; // @[addsub_64.scala 39:22]
  assign fa_12_io_i0 = io_i0[12]; // @[addsub_64.scala 37:29]
  assign fa_12_io_i1 = io_onesComp_ip[12]; // @[addsub_64.scala 38:38]
  assign fa_12_io_cin = fa_11_io_cout; // @[addsub_64.scala 39:22]
  assign fa_13_io_i0 = io_i0[13]; // @[addsub_64.scala 37:29]
  assign fa_13_io_i1 = io_onesComp_ip[13]; // @[addsub_64.scala 38:38]
  assign fa_13_io_cin = fa_12_io_cout; // @[addsub_64.scala 39:22]
  assign fa_14_io_i0 = io_i0[14]; // @[addsub_64.scala 37:29]
  assign fa_14_io_i1 = io_onesComp_ip[14]; // @[addsub_64.scala 38:38]
  assign fa_14_io_cin = fa_13_io_cout; // @[addsub_64.scala 39:22]
  assign fa_15_io_i0 = io_i0[15]; // @[addsub_64.scala 37:29]
  assign fa_15_io_i1 = io_onesComp_ip[15]; // @[addsub_64.scala 38:38]
  assign fa_15_io_cin = fa_14_io_cout; // @[addsub_64.scala 39:22]
  assign fa_16_io_i0 = io_i0[16]; // @[addsub_64.scala 37:29]
  assign fa_16_io_i1 = io_onesComp_ip[16]; // @[addsub_64.scala 38:38]
  assign fa_16_io_cin = fa_15_io_cout; // @[addsub_64.scala 39:22]
  assign fa_17_io_i0 = io_i0[17]; // @[addsub_64.scala 37:29]
  assign fa_17_io_i1 = io_onesComp_ip[17]; // @[addsub_64.scala 38:38]
  assign fa_17_io_cin = fa_16_io_cout; // @[addsub_64.scala 39:22]
  assign fa_18_io_i0 = io_i0[18]; // @[addsub_64.scala 37:29]
  assign fa_18_io_i1 = io_onesComp_ip[18]; // @[addsub_64.scala 38:38]
  assign fa_18_io_cin = fa_17_io_cout; // @[addsub_64.scala 39:22]
  assign fa_19_io_i0 = io_i0[19]; // @[addsub_64.scala 37:29]
  assign fa_19_io_i1 = io_onesComp_ip[19]; // @[addsub_64.scala 38:38]
  assign fa_19_io_cin = fa_18_io_cout; // @[addsub_64.scala 39:22]
  assign fa_20_io_i0 = io_i0[20]; // @[addsub_64.scala 37:29]
  assign fa_20_io_i1 = io_onesComp_ip[20]; // @[addsub_64.scala 38:38]
  assign fa_20_io_cin = fa_19_io_cout; // @[addsub_64.scala 39:22]
  assign fa_21_io_i0 = io_i0[21]; // @[addsub_64.scala 37:29]
  assign fa_21_io_i1 = io_onesComp_ip[21]; // @[addsub_64.scala 38:38]
  assign fa_21_io_cin = fa_20_io_cout; // @[addsub_64.scala 39:22]
  assign fa_22_io_i0 = io_i0[22]; // @[addsub_64.scala 37:29]
  assign fa_22_io_i1 = io_onesComp_ip[22]; // @[addsub_64.scala 38:38]
  assign fa_22_io_cin = fa_21_io_cout; // @[addsub_64.scala 39:22]
  assign fa_23_io_i0 = io_i0[23]; // @[addsub_64.scala 37:29]
  assign fa_23_io_i1 = io_onesComp_ip[23]; // @[addsub_64.scala 38:38]
  assign fa_23_io_cin = fa_22_io_cout; // @[addsub_64.scala 39:22]
  assign fa_24_io_i0 = io_i0[24]; // @[addsub_64.scala 37:29]
  assign fa_24_io_i1 = io_onesComp_ip[24]; // @[addsub_64.scala 38:38]
  assign fa_24_io_cin = fa_23_io_cout; // @[addsub_64.scala 39:22]
  assign fa_25_io_i0 = io_i0[25]; // @[addsub_64.scala 37:29]
  assign fa_25_io_i1 = io_onesComp_ip[25]; // @[addsub_64.scala 38:38]
  assign fa_25_io_cin = fa_24_io_cout; // @[addsub_64.scala 39:22]
  assign fa_26_io_i0 = io_i0[26]; // @[addsub_64.scala 37:29]
  assign fa_26_io_i1 = io_onesComp_ip[26]; // @[addsub_64.scala 38:38]
  assign fa_26_io_cin = fa_25_io_cout; // @[addsub_64.scala 39:22]
  assign fa_27_io_i0 = io_i0[27]; // @[addsub_64.scala 37:29]
  assign fa_27_io_i1 = io_onesComp_ip[27]; // @[addsub_64.scala 38:38]
  assign fa_27_io_cin = fa_26_io_cout; // @[addsub_64.scala 39:22]
  assign fa_28_io_i0 = io_i0[28]; // @[addsub_64.scala 37:29]
  assign fa_28_io_i1 = io_onesComp_ip[28]; // @[addsub_64.scala 38:38]
  assign fa_28_io_cin = fa_27_io_cout; // @[addsub_64.scala 39:22]
  assign fa_29_io_i0 = io_i0[29]; // @[addsub_64.scala 37:29]
  assign fa_29_io_i1 = io_onesComp_ip[29]; // @[addsub_64.scala 38:38]
  assign fa_29_io_cin = fa_28_io_cout; // @[addsub_64.scala 39:22]
  assign fa_30_io_i0 = io_i0[30]; // @[addsub_64.scala 37:29]
  assign fa_30_io_i1 = io_onesComp_ip[30]; // @[addsub_64.scala 38:38]
  assign fa_30_io_cin = fa_29_io_cout; // @[addsub_64.scala 39:22]
  assign fa_31_io_i0 = io_i0[31]; // @[addsub_64.scala 37:29]
  assign fa_31_io_i1 = io_onesComp_ip[31]; // @[addsub_64.scala 38:38]
  assign fa_31_io_cin = fa_30_io_cout; // @[addsub_64.scala 39:22]
  assign fa_32_io_i0 = io_i0[32]; // @[addsub_64.scala 37:29]
  assign fa_32_io_i1 = io_onesComp_ip[32]; // @[addsub_64.scala 38:38]
  assign fa_32_io_cin = fa_31_io_cout; // @[addsub_64.scala 39:22]
  assign fa_33_io_i0 = io_i0[33]; // @[addsub_64.scala 37:29]
  assign fa_33_io_i1 = io_onesComp_ip[33]; // @[addsub_64.scala 38:38]
  assign fa_33_io_cin = fa_32_io_cout; // @[addsub_64.scala 39:22]
  assign fa_34_io_i0 = io_i0[34]; // @[addsub_64.scala 37:29]
  assign fa_34_io_i1 = io_onesComp_ip[34]; // @[addsub_64.scala 38:38]
  assign fa_34_io_cin = fa_33_io_cout; // @[addsub_64.scala 39:22]
  assign fa_35_io_i0 = io_i0[35]; // @[addsub_64.scala 37:29]
  assign fa_35_io_i1 = io_onesComp_ip[35]; // @[addsub_64.scala 38:38]
  assign fa_35_io_cin = fa_34_io_cout; // @[addsub_64.scala 39:22]
  assign fa_36_io_i0 = io_i0[36]; // @[addsub_64.scala 37:29]
  assign fa_36_io_i1 = io_onesComp_ip[36]; // @[addsub_64.scala 38:38]
  assign fa_36_io_cin = fa_35_io_cout; // @[addsub_64.scala 39:22]
  assign fa_37_io_i0 = io_i0[37]; // @[addsub_64.scala 37:29]
  assign fa_37_io_i1 = io_onesComp_ip[37]; // @[addsub_64.scala 38:38]
  assign fa_37_io_cin = fa_36_io_cout; // @[addsub_64.scala 39:22]
  assign fa_38_io_i0 = io_i0[38]; // @[addsub_64.scala 37:29]
  assign fa_38_io_i1 = io_onesComp_ip[38]; // @[addsub_64.scala 38:38]
  assign fa_38_io_cin = fa_37_io_cout; // @[addsub_64.scala 39:22]
  assign fa_39_io_i0 = io_i0[39]; // @[addsub_64.scala 37:29]
  assign fa_39_io_i1 = io_onesComp_ip[39]; // @[addsub_64.scala 38:38]
  assign fa_39_io_cin = fa_38_io_cout; // @[addsub_64.scala 39:22]
  assign fa_40_io_i0 = io_i0[40]; // @[addsub_64.scala 37:29]
  assign fa_40_io_i1 = io_onesComp_ip[40]; // @[addsub_64.scala 38:38]
  assign fa_40_io_cin = fa_39_io_cout; // @[addsub_64.scala 39:22]
  assign fa_41_io_i0 = io_i0[41]; // @[addsub_64.scala 37:29]
  assign fa_41_io_i1 = io_onesComp_ip[41]; // @[addsub_64.scala 38:38]
  assign fa_41_io_cin = fa_40_io_cout; // @[addsub_64.scala 39:22]
  assign fa_42_io_i0 = io_i0[42]; // @[addsub_64.scala 37:29]
  assign fa_42_io_i1 = io_onesComp_ip[42]; // @[addsub_64.scala 38:38]
  assign fa_42_io_cin = fa_41_io_cout; // @[addsub_64.scala 39:22]
  assign fa_43_io_i0 = io_i0[43]; // @[addsub_64.scala 37:29]
  assign fa_43_io_i1 = io_onesComp_ip[43]; // @[addsub_64.scala 38:38]
  assign fa_43_io_cin = fa_42_io_cout; // @[addsub_64.scala 39:22]
  assign fa_44_io_i0 = io_i0[44]; // @[addsub_64.scala 37:29]
  assign fa_44_io_i1 = io_onesComp_ip[44]; // @[addsub_64.scala 38:38]
  assign fa_44_io_cin = fa_43_io_cout; // @[addsub_64.scala 39:22]
  assign fa_45_io_i0 = io_i0[45]; // @[addsub_64.scala 37:29]
  assign fa_45_io_i1 = io_onesComp_ip[45]; // @[addsub_64.scala 38:38]
  assign fa_45_io_cin = fa_44_io_cout; // @[addsub_64.scala 39:22]
  assign fa_46_io_i0 = io_i0[46]; // @[addsub_64.scala 37:29]
  assign fa_46_io_i1 = io_onesComp_ip[46]; // @[addsub_64.scala 38:38]
  assign fa_46_io_cin = fa_45_io_cout; // @[addsub_64.scala 39:22]
  assign fa_47_io_i0 = io_i0[47]; // @[addsub_64.scala 37:29]
  assign fa_47_io_i1 = io_onesComp_ip[47]; // @[addsub_64.scala 38:38]
  assign fa_47_io_cin = fa_46_io_cout; // @[addsub_64.scala 39:22]
  assign fa_48_io_i0 = io_i0[48]; // @[addsub_64.scala 37:29]
  assign fa_48_io_i1 = io_onesComp_ip[48]; // @[addsub_64.scala 38:38]
  assign fa_48_io_cin = fa_47_io_cout; // @[addsub_64.scala 39:22]
  assign fa_49_io_i0 = io_i0[49]; // @[addsub_64.scala 37:29]
  assign fa_49_io_i1 = io_onesComp_ip[49]; // @[addsub_64.scala 38:38]
  assign fa_49_io_cin = fa_48_io_cout; // @[addsub_64.scala 39:22]
  assign fa_50_io_i0 = io_i0[50]; // @[addsub_64.scala 37:29]
  assign fa_50_io_i1 = io_onesComp_ip[50]; // @[addsub_64.scala 38:38]
  assign fa_50_io_cin = fa_49_io_cout; // @[addsub_64.scala 39:22]
  assign fa_51_io_i0 = io_i0[51]; // @[addsub_64.scala 37:29]
  assign fa_51_io_i1 = io_onesComp_ip[51]; // @[addsub_64.scala 38:38]
  assign fa_51_io_cin = fa_50_io_cout; // @[addsub_64.scala 39:22]
  assign fa_52_io_i0 = io_i0[52]; // @[addsub_64.scala 37:29]
  assign fa_52_io_i1 = io_onesComp_ip[52]; // @[addsub_64.scala 38:38]
  assign fa_52_io_cin = fa_51_io_cout; // @[addsub_64.scala 39:22]
  assign fa_53_io_i0 = io_i0[53]; // @[addsub_64.scala 37:29]
  assign fa_53_io_i1 = io_onesComp_ip[53]; // @[addsub_64.scala 38:38]
  assign fa_53_io_cin = fa_52_io_cout; // @[addsub_64.scala 39:22]
  assign fa_54_io_i0 = io_i0[54]; // @[addsub_64.scala 37:29]
  assign fa_54_io_i1 = io_onesComp_ip[54]; // @[addsub_64.scala 38:38]
  assign fa_54_io_cin = fa_53_io_cout; // @[addsub_64.scala 39:22]
  assign fa_55_io_i0 = io_i0[55]; // @[addsub_64.scala 37:29]
  assign fa_55_io_i1 = io_onesComp_ip[55]; // @[addsub_64.scala 38:38]
  assign fa_55_io_cin = fa_54_io_cout; // @[addsub_64.scala 39:22]
  assign fa_56_io_i0 = io_i0[56]; // @[addsub_64.scala 37:29]
  assign fa_56_io_i1 = io_onesComp_ip[56]; // @[addsub_64.scala 38:38]
  assign fa_56_io_cin = fa_55_io_cout; // @[addsub_64.scala 39:22]
  assign fa_57_io_i0 = io_i0[57]; // @[addsub_64.scala 37:29]
  assign fa_57_io_i1 = io_onesComp_ip[57]; // @[addsub_64.scala 38:38]
  assign fa_57_io_cin = fa_56_io_cout; // @[addsub_64.scala 39:22]
  assign fa_58_io_i0 = io_i0[58]; // @[addsub_64.scala 37:29]
  assign fa_58_io_i1 = io_onesComp_ip[58]; // @[addsub_64.scala 38:38]
  assign fa_58_io_cin = fa_57_io_cout; // @[addsub_64.scala 39:22]
  assign fa_59_io_i0 = io_i0[59]; // @[addsub_64.scala 37:29]
  assign fa_59_io_i1 = io_onesComp_ip[59]; // @[addsub_64.scala 38:38]
  assign fa_59_io_cin = fa_58_io_cout; // @[addsub_64.scala 39:22]
  assign fa_60_io_i0 = io_i0[60]; // @[addsub_64.scala 37:29]
  assign fa_60_io_i1 = io_onesComp_ip[60]; // @[addsub_64.scala 38:38]
  assign fa_60_io_cin = fa_59_io_cout; // @[addsub_64.scala 39:22]
  assign fa_61_io_i0 = io_i0[61]; // @[addsub_64.scala 37:29]
  assign fa_61_io_i1 = io_onesComp_ip[61]; // @[addsub_64.scala 38:38]
  assign fa_61_io_cin = fa_60_io_cout; // @[addsub_64.scala 39:22]
  assign fa_62_io_i0 = io_i0[62]; // @[addsub_64.scala 37:29]
  assign fa_62_io_i1 = io_onesComp_ip[62]; // @[addsub_64.scala 38:38]
  assign fa_62_io_cin = fa_61_io_cout; // @[addsub_64.scala 39:22]
  assign fa_63_io_i0 = io_i0[63]; // @[addsub_64.scala 37:29]
  assign fa_63_io_i1 = io_onesComp_ip[63]; // @[addsub_64.scala 38:38]
  assign fa_63_io_cin = fa_62_io_cout; // @[addsub_64.scala 39:22]
endmodule
