module xor2(
  input   io_a,
  output  io_out
);
  assign io_out = io_a ^ 1'h1; // @[getOnesComplement.scala 13:20]
endmodule
module getOnesComplement(
  input  [63:0] io_i1,
  output [63:0] io_onesComp
);
  wire  xor_0_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_0_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_1_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_1_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_2_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_2_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_3_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_3_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_4_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_4_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_5_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_5_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_6_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_6_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_7_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_7_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_8_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_8_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_9_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_9_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_10_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_10_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_11_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_11_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_12_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_12_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_13_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_13_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_14_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_14_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_15_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_15_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_16_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_16_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_17_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_17_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_18_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_18_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_19_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_19_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_20_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_20_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_21_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_21_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_22_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_22_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_23_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_23_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_24_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_24_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_25_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_25_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_26_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_26_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_27_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_27_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_28_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_28_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_29_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_29_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_30_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_30_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_31_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_31_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_32_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_32_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_33_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_33_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_34_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_34_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_35_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_35_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_36_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_36_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_37_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_37_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_38_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_38_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_39_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_39_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_40_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_40_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_41_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_41_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_42_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_42_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_43_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_43_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_44_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_44_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_45_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_45_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_46_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_46_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_47_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_47_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_48_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_48_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_49_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_49_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_50_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_50_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_51_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_51_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_52_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_52_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_53_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_53_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_54_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_54_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_55_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_55_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_56_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_56_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_57_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_57_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_58_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_58_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_59_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_59_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_60_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_60_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_61_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_61_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_62_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_62_io_out; // @[getOnesComplement.scala 24:33]
  wire  xor_63_io_a; // @[getOnesComplement.scala 24:33]
  wire  xor_63_io_out; // @[getOnesComplement.scala 24:33]
  wire [7:0] lo_lo_lo = {xor_7_io_out,xor_6_io_out,xor_5_io_out,xor_4_io_out,xor_3_io_out,xor_2_io_out,xor_1_io_out,
    xor_0_io_out}; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {xor_15_io_out,xor_14_io_out,xor_13_io_out,xor_12_io_out,xor_11_io_out,xor_10_io_out,xor_9_io_out,
    xor_8_io_out,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {xor_23_io_out,xor_22_io_out,xor_21_io_out,xor_20_io_out,xor_19_io_out,xor_18_io_out,
    xor_17_io_out,xor_16_io_out}; // @[Cat.scala 30:58]
  wire [31:0] lo = {xor_31_io_out,xor_30_io_out,xor_29_io_out,xor_28_io_out,xor_27_io_out,xor_26_io_out,xor_25_io_out,
    xor_24_io_out,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {xor_39_io_out,xor_38_io_out,xor_37_io_out,xor_36_io_out,xor_35_io_out,xor_34_io_out,
    xor_33_io_out,xor_32_io_out}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {xor_47_io_out,xor_46_io_out,xor_45_io_out,xor_44_io_out,xor_43_io_out,xor_42_io_out,xor_41_io_out
    ,xor_40_io_out,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {xor_55_io_out,xor_54_io_out,xor_53_io_out,xor_52_io_out,xor_51_io_out,xor_50_io_out,
    xor_49_io_out,xor_48_io_out}; // @[Cat.scala 30:58]
  wire [31:0] hi = {xor_63_io_out,xor_62_io_out,xor_61_io_out,xor_60_io_out,xor_59_io_out,xor_58_io_out,xor_57_io_out,
    xor_56_io_out,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  xor2 xor_0 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_0_io_a),
    .io_out(xor_0_io_out)
  );
  xor2 xor_1 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_1_io_a),
    .io_out(xor_1_io_out)
  );
  xor2 xor_2 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_2_io_a),
    .io_out(xor_2_io_out)
  );
  xor2 xor_3 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_3_io_a),
    .io_out(xor_3_io_out)
  );
  xor2 xor_4 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_4_io_a),
    .io_out(xor_4_io_out)
  );
  xor2 xor_5 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_5_io_a),
    .io_out(xor_5_io_out)
  );
  xor2 xor_6 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_6_io_a),
    .io_out(xor_6_io_out)
  );
  xor2 xor_7 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_7_io_a),
    .io_out(xor_7_io_out)
  );
  xor2 xor_8 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_8_io_a),
    .io_out(xor_8_io_out)
  );
  xor2 xor_9 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_9_io_a),
    .io_out(xor_9_io_out)
  );
  xor2 xor_10 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_10_io_a),
    .io_out(xor_10_io_out)
  );
  xor2 xor_11 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_11_io_a),
    .io_out(xor_11_io_out)
  );
  xor2 xor_12 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_12_io_a),
    .io_out(xor_12_io_out)
  );
  xor2 xor_13 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_13_io_a),
    .io_out(xor_13_io_out)
  );
  xor2 xor_14 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_14_io_a),
    .io_out(xor_14_io_out)
  );
  xor2 xor_15 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_15_io_a),
    .io_out(xor_15_io_out)
  );
  xor2 xor_16 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_16_io_a),
    .io_out(xor_16_io_out)
  );
  xor2 xor_17 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_17_io_a),
    .io_out(xor_17_io_out)
  );
  xor2 xor_18 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_18_io_a),
    .io_out(xor_18_io_out)
  );
  xor2 xor_19 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_19_io_a),
    .io_out(xor_19_io_out)
  );
  xor2 xor_20 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_20_io_a),
    .io_out(xor_20_io_out)
  );
  xor2 xor_21 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_21_io_a),
    .io_out(xor_21_io_out)
  );
  xor2 xor_22 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_22_io_a),
    .io_out(xor_22_io_out)
  );
  xor2 xor_23 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_23_io_a),
    .io_out(xor_23_io_out)
  );
  xor2 xor_24 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_24_io_a),
    .io_out(xor_24_io_out)
  );
  xor2 xor_25 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_25_io_a),
    .io_out(xor_25_io_out)
  );
  xor2 xor_26 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_26_io_a),
    .io_out(xor_26_io_out)
  );
  xor2 xor_27 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_27_io_a),
    .io_out(xor_27_io_out)
  );
  xor2 xor_28 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_28_io_a),
    .io_out(xor_28_io_out)
  );
  xor2 xor_29 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_29_io_a),
    .io_out(xor_29_io_out)
  );
  xor2 xor_30 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_30_io_a),
    .io_out(xor_30_io_out)
  );
  xor2 xor_31 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_31_io_a),
    .io_out(xor_31_io_out)
  );
  xor2 xor_32 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_32_io_a),
    .io_out(xor_32_io_out)
  );
  xor2 xor_33 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_33_io_a),
    .io_out(xor_33_io_out)
  );
  xor2 xor_34 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_34_io_a),
    .io_out(xor_34_io_out)
  );
  xor2 xor_35 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_35_io_a),
    .io_out(xor_35_io_out)
  );
  xor2 xor_36 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_36_io_a),
    .io_out(xor_36_io_out)
  );
  xor2 xor_37 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_37_io_a),
    .io_out(xor_37_io_out)
  );
  xor2 xor_38 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_38_io_a),
    .io_out(xor_38_io_out)
  );
  xor2 xor_39 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_39_io_a),
    .io_out(xor_39_io_out)
  );
  xor2 xor_40 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_40_io_a),
    .io_out(xor_40_io_out)
  );
  xor2 xor_41 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_41_io_a),
    .io_out(xor_41_io_out)
  );
  xor2 xor_42 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_42_io_a),
    .io_out(xor_42_io_out)
  );
  xor2 xor_43 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_43_io_a),
    .io_out(xor_43_io_out)
  );
  xor2 xor_44 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_44_io_a),
    .io_out(xor_44_io_out)
  );
  xor2 xor_45 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_45_io_a),
    .io_out(xor_45_io_out)
  );
  xor2 xor_46 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_46_io_a),
    .io_out(xor_46_io_out)
  );
  xor2 xor_47 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_47_io_a),
    .io_out(xor_47_io_out)
  );
  xor2 xor_48 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_48_io_a),
    .io_out(xor_48_io_out)
  );
  xor2 xor_49 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_49_io_a),
    .io_out(xor_49_io_out)
  );
  xor2 xor_50 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_50_io_a),
    .io_out(xor_50_io_out)
  );
  xor2 xor_51 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_51_io_a),
    .io_out(xor_51_io_out)
  );
  xor2 xor_52 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_52_io_a),
    .io_out(xor_52_io_out)
  );
  xor2 xor_53 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_53_io_a),
    .io_out(xor_53_io_out)
  );
  xor2 xor_54 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_54_io_a),
    .io_out(xor_54_io_out)
  );
  xor2 xor_55 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_55_io_a),
    .io_out(xor_55_io_out)
  );
  xor2 xor_56 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_56_io_a),
    .io_out(xor_56_io_out)
  );
  xor2 xor_57 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_57_io_a),
    .io_out(xor_57_io_out)
  );
  xor2 xor_58 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_58_io_a),
    .io_out(xor_58_io_out)
  );
  xor2 xor_59 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_59_io_a),
    .io_out(xor_59_io_out)
  );
  xor2 xor_60 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_60_io_a),
    .io_out(xor_60_io_out)
  );
  xor2 xor_61 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_61_io_a),
    .io_out(xor_61_io_out)
  );
  xor2 xor_62 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_62_io_a),
    .io_out(xor_62_io_out)
  );
  xor2 xor_63 ( // @[getOnesComplement.scala 24:33]
    .io_a(xor_63_io_a),
    .io_out(xor_63_io_out)
  );
  assign io_onesComp = {hi,lo}; // @[Cat.scala 30:58]
  assign xor_0_io_a = io_i1[0]; // @[getOnesComplement.scala 27:29]
  assign xor_1_io_a = io_i1[1]; // @[getOnesComplement.scala 27:29]
  assign xor_2_io_a = io_i1[2]; // @[getOnesComplement.scala 27:29]
  assign xor_3_io_a = io_i1[3]; // @[getOnesComplement.scala 27:29]
  assign xor_4_io_a = io_i1[4]; // @[getOnesComplement.scala 27:29]
  assign xor_5_io_a = io_i1[5]; // @[getOnesComplement.scala 27:29]
  assign xor_6_io_a = io_i1[6]; // @[getOnesComplement.scala 27:29]
  assign xor_7_io_a = io_i1[7]; // @[getOnesComplement.scala 27:29]
  assign xor_8_io_a = io_i1[8]; // @[getOnesComplement.scala 27:29]
  assign xor_9_io_a = io_i1[9]; // @[getOnesComplement.scala 27:29]
  assign xor_10_io_a = io_i1[10]; // @[getOnesComplement.scala 27:29]
  assign xor_11_io_a = io_i1[11]; // @[getOnesComplement.scala 27:29]
  assign xor_12_io_a = io_i1[12]; // @[getOnesComplement.scala 27:29]
  assign xor_13_io_a = io_i1[13]; // @[getOnesComplement.scala 27:29]
  assign xor_14_io_a = io_i1[14]; // @[getOnesComplement.scala 27:29]
  assign xor_15_io_a = io_i1[15]; // @[getOnesComplement.scala 27:29]
  assign xor_16_io_a = io_i1[16]; // @[getOnesComplement.scala 27:29]
  assign xor_17_io_a = io_i1[17]; // @[getOnesComplement.scala 27:29]
  assign xor_18_io_a = io_i1[18]; // @[getOnesComplement.scala 27:29]
  assign xor_19_io_a = io_i1[19]; // @[getOnesComplement.scala 27:29]
  assign xor_20_io_a = io_i1[20]; // @[getOnesComplement.scala 27:29]
  assign xor_21_io_a = io_i1[21]; // @[getOnesComplement.scala 27:29]
  assign xor_22_io_a = io_i1[22]; // @[getOnesComplement.scala 27:29]
  assign xor_23_io_a = io_i1[23]; // @[getOnesComplement.scala 27:29]
  assign xor_24_io_a = io_i1[24]; // @[getOnesComplement.scala 27:29]
  assign xor_25_io_a = io_i1[25]; // @[getOnesComplement.scala 27:29]
  assign xor_26_io_a = io_i1[26]; // @[getOnesComplement.scala 27:29]
  assign xor_27_io_a = io_i1[27]; // @[getOnesComplement.scala 27:29]
  assign xor_28_io_a = io_i1[28]; // @[getOnesComplement.scala 27:29]
  assign xor_29_io_a = io_i1[29]; // @[getOnesComplement.scala 27:29]
  assign xor_30_io_a = io_i1[30]; // @[getOnesComplement.scala 27:29]
  assign xor_31_io_a = io_i1[31]; // @[getOnesComplement.scala 27:29]
  assign xor_32_io_a = io_i1[32]; // @[getOnesComplement.scala 27:29]
  assign xor_33_io_a = io_i1[33]; // @[getOnesComplement.scala 27:29]
  assign xor_34_io_a = io_i1[34]; // @[getOnesComplement.scala 27:29]
  assign xor_35_io_a = io_i1[35]; // @[getOnesComplement.scala 27:29]
  assign xor_36_io_a = io_i1[36]; // @[getOnesComplement.scala 27:29]
  assign xor_37_io_a = io_i1[37]; // @[getOnesComplement.scala 27:29]
  assign xor_38_io_a = io_i1[38]; // @[getOnesComplement.scala 27:29]
  assign xor_39_io_a = io_i1[39]; // @[getOnesComplement.scala 27:29]
  assign xor_40_io_a = io_i1[40]; // @[getOnesComplement.scala 27:29]
  assign xor_41_io_a = io_i1[41]; // @[getOnesComplement.scala 27:29]
  assign xor_42_io_a = io_i1[42]; // @[getOnesComplement.scala 27:29]
  assign xor_43_io_a = io_i1[43]; // @[getOnesComplement.scala 27:29]
  assign xor_44_io_a = io_i1[44]; // @[getOnesComplement.scala 27:29]
  assign xor_45_io_a = io_i1[45]; // @[getOnesComplement.scala 27:29]
  assign xor_46_io_a = io_i1[46]; // @[getOnesComplement.scala 27:29]
  assign xor_47_io_a = io_i1[47]; // @[getOnesComplement.scala 27:29]
  assign xor_48_io_a = io_i1[48]; // @[getOnesComplement.scala 27:29]
  assign xor_49_io_a = io_i1[49]; // @[getOnesComplement.scala 27:29]
  assign xor_50_io_a = io_i1[50]; // @[getOnesComplement.scala 27:29]
  assign xor_51_io_a = io_i1[51]; // @[getOnesComplement.scala 27:29]
  assign xor_52_io_a = io_i1[52]; // @[getOnesComplement.scala 27:29]
  assign xor_53_io_a = io_i1[53]; // @[getOnesComplement.scala 27:29]
  assign xor_54_io_a = io_i1[54]; // @[getOnesComplement.scala 27:29]
  assign xor_55_io_a = io_i1[55]; // @[getOnesComplement.scala 27:29]
  assign xor_56_io_a = io_i1[56]; // @[getOnesComplement.scala 27:29]
  assign xor_57_io_a = io_i1[57]; // @[getOnesComplement.scala 27:29]
  assign xor_58_io_a = io_i1[58]; // @[getOnesComplement.scala 27:29]
  assign xor_59_io_a = io_i1[59]; // @[getOnesComplement.scala 27:29]
  assign xor_60_io_a = io_i1[60]; // @[getOnesComplement.scala 27:29]
  assign xor_61_io_a = io_i1[61]; // @[getOnesComplement.scala 27:29]
  assign xor_62_io_a = io_i1[62]; // @[getOnesComplement.scala 27:29]
  assign xor_63_io_a = io_i1[63]; // @[getOnesComplement.scala 27:29]
endmodule
module fullAdder(
  input   io_i0,
  input   io_i1,
  input   io_cin,
  output  io_sum,
  output  io_cout
);
  assign io_sum = io_i0 ^ io_i1 ^ io_cin; // @[addsub.scala 14:29]
  assign io_cout = io_i0 & io_i1 | io_i1 & io_cin | io_cin & io_i0; // @[addsub.scala 15:51]
endmodule
module addsub(
  input  [63:0] io_onesComp_ip,
  input  [63:0] io_i0,
  output [63:0] io_sum
);
  wire  fa_0_io_i0; // @[addsub.scala 28:32]
  wire  fa_0_io_i1; // @[addsub.scala 28:32]
  wire  fa_0_io_cin; // @[addsub.scala 28:32]
  wire  fa_0_io_sum; // @[addsub.scala 28:32]
  wire  fa_0_io_cout; // @[addsub.scala 28:32]
  wire  fa_1_io_i0; // @[addsub.scala 28:32]
  wire  fa_1_io_i1; // @[addsub.scala 28:32]
  wire  fa_1_io_cin; // @[addsub.scala 28:32]
  wire  fa_1_io_sum; // @[addsub.scala 28:32]
  wire  fa_1_io_cout; // @[addsub.scala 28:32]
  wire  fa_2_io_i0; // @[addsub.scala 28:32]
  wire  fa_2_io_i1; // @[addsub.scala 28:32]
  wire  fa_2_io_cin; // @[addsub.scala 28:32]
  wire  fa_2_io_sum; // @[addsub.scala 28:32]
  wire  fa_2_io_cout; // @[addsub.scala 28:32]
  wire  fa_3_io_i0; // @[addsub.scala 28:32]
  wire  fa_3_io_i1; // @[addsub.scala 28:32]
  wire  fa_3_io_cin; // @[addsub.scala 28:32]
  wire  fa_3_io_sum; // @[addsub.scala 28:32]
  wire  fa_3_io_cout; // @[addsub.scala 28:32]
  wire  fa_4_io_i0; // @[addsub.scala 28:32]
  wire  fa_4_io_i1; // @[addsub.scala 28:32]
  wire  fa_4_io_cin; // @[addsub.scala 28:32]
  wire  fa_4_io_sum; // @[addsub.scala 28:32]
  wire  fa_4_io_cout; // @[addsub.scala 28:32]
  wire  fa_5_io_i0; // @[addsub.scala 28:32]
  wire  fa_5_io_i1; // @[addsub.scala 28:32]
  wire  fa_5_io_cin; // @[addsub.scala 28:32]
  wire  fa_5_io_sum; // @[addsub.scala 28:32]
  wire  fa_5_io_cout; // @[addsub.scala 28:32]
  wire  fa_6_io_i0; // @[addsub.scala 28:32]
  wire  fa_6_io_i1; // @[addsub.scala 28:32]
  wire  fa_6_io_cin; // @[addsub.scala 28:32]
  wire  fa_6_io_sum; // @[addsub.scala 28:32]
  wire  fa_6_io_cout; // @[addsub.scala 28:32]
  wire  fa_7_io_i0; // @[addsub.scala 28:32]
  wire  fa_7_io_i1; // @[addsub.scala 28:32]
  wire  fa_7_io_cin; // @[addsub.scala 28:32]
  wire  fa_7_io_sum; // @[addsub.scala 28:32]
  wire  fa_7_io_cout; // @[addsub.scala 28:32]
  wire  fa_8_io_i0; // @[addsub.scala 28:32]
  wire  fa_8_io_i1; // @[addsub.scala 28:32]
  wire  fa_8_io_cin; // @[addsub.scala 28:32]
  wire  fa_8_io_sum; // @[addsub.scala 28:32]
  wire  fa_8_io_cout; // @[addsub.scala 28:32]
  wire  fa_9_io_i0; // @[addsub.scala 28:32]
  wire  fa_9_io_i1; // @[addsub.scala 28:32]
  wire  fa_9_io_cin; // @[addsub.scala 28:32]
  wire  fa_9_io_sum; // @[addsub.scala 28:32]
  wire  fa_9_io_cout; // @[addsub.scala 28:32]
  wire  fa_10_io_i0; // @[addsub.scala 28:32]
  wire  fa_10_io_i1; // @[addsub.scala 28:32]
  wire  fa_10_io_cin; // @[addsub.scala 28:32]
  wire  fa_10_io_sum; // @[addsub.scala 28:32]
  wire  fa_10_io_cout; // @[addsub.scala 28:32]
  wire  fa_11_io_i0; // @[addsub.scala 28:32]
  wire  fa_11_io_i1; // @[addsub.scala 28:32]
  wire  fa_11_io_cin; // @[addsub.scala 28:32]
  wire  fa_11_io_sum; // @[addsub.scala 28:32]
  wire  fa_11_io_cout; // @[addsub.scala 28:32]
  wire  fa_12_io_i0; // @[addsub.scala 28:32]
  wire  fa_12_io_i1; // @[addsub.scala 28:32]
  wire  fa_12_io_cin; // @[addsub.scala 28:32]
  wire  fa_12_io_sum; // @[addsub.scala 28:32]
  wire  fa_12_io_cout; // @[addsub.scala 28:32]
  wire  fa_13_io_i0; // @[addsub.scala 28:32]
  wire  fa_13_io_i1; // @[addsub.scala 28:32]
  wire  fa_13_io_cin; // @[addsub.scala 28:32]
  wire  fa_13_io_sum; // @[addsub.scala 28:32]
  wire  fa_13_io_cout; // @[addsub.scala 28:32]
  wire  fa_14_io_i0; // @[addsub.scala 28:32]
  wire  fa_14_io_i1; // @[addsub.scala 28:32]
  wire  fa_14_io_cin; // @[addsub.scala 28:32]
  wire  fa_14_io_sum; // @[addsub.scala 28:32]
  wire  fa_14_io_cout; // @[addsub.scala 28:32]
  wire  fa_15_io_i0; // @[addsub.scala 28:32]
  wire  fa_15_io_i1; // @[addsub.scala 28:32]
  wire  fa_15_io_cin; // @[addsub.scala 28:32]
  wire  fa_15_io_sum; // @[addsub.scala 28:32]
  wire  fa_15_io_cout; // @[addsub.scala 28:32]
  wire  fa_16_io_i0; // @[addsub.scala 28:32]
  wire  fa_16_io_i1; // @[addsub.scala 28:32]
  wire  fa_16_io_cin; // @[addsub.scala 28:32]
  wire  fa_16_io_sum; // @[addsub.scala 28:32]
  wire  fa_16_io_cout; // @[addsub.scala 28:32]
  wire  fa_17_io_i0; // @[addsub.scala 28:32]
  wire  fa_17_io_i1; // @[addsub.scala 28:32]
  wire  fa_17_io_cin; // @[addsub.scala 28:32]
  wire  fa_17_io_sum; // @[addsub.scala 28:32]
  wire  fa_17_io_cout; // @[addsub.scala 28:32]
  wire  fa_18_io_i0; // @[addsub.scala 28:32]
  wire  fa_18_io_i1; // @[addsub.scala 28:32]
  wire  fa_18_io_cin; // @[addsub.scala 28:32]
  wire  fa_18_io_sum; // @[addsub.scala 28:32]
  wire  fa_18_io_cout; // @[addsub.scala 28:32]
  wire  fa_19_io_i0; // @[addsub.scala 28:32]
  wire  fa_19_io_i1; // @[addsub.scala 28:32]
  wire  fa_19_io_cin; // @[addsub.scala 28:32]
  wire  fa_19_io_sum; // @[addsub.scala 28:32]
  wire  fa_19_io_cout; // @[addsub.scala 28:32]
  wire  fa_20_io_i0; // @[addsub.scala 28:32]
  wire  fa_20_io_i1; // @[addsub.scala 28:32]
  wire  fa_20_io_cin; // @[addsub.scala 28:32]
  wire  fa_20_io_sum; // @[addsub.scala 28:32]
  wire  fa_20_io_cout; // @[addsub.scala 28:32]
  wire  fa_21_io_i0; // @[addsub.scala 28:32]
  wire  fa_21_io_i1; // @[addsub.scala 28:32]
  wire  fa_21_io_cin; // @[addsub.scala 28:32]
  wire  fa_21_io_sum; // @[addsub.scala 28:32]
  wire  fa_21_io_cout; // @[addsub.scala 28:32]
  wire  fa_22_io_i0; // @[addsub.scala 28:32]
  wire  fa_22_io_i1; // @[addsub.scala 28:32]
  wire  fa_22_io_cin; // @[addsub.scala 28:32]
  wire  fa_22_io_sum; // @[addsub.scala 28:32]
  wire  fa_22_io_cout; // @[addsub.scala 28:32]
  wire  fa_23_io_i0; // @[addsub.scala 28:32]
  wire  fa_23_io_i1; // @[addsub.scala 28:32]
  wire  fa_23_io_cin; // @[addsub.scala 28:32]
  wire  fa_23_io_sum; // @[addsub.scala 28:32]
  wire  fa_23_io_cout; // @[addsub.scala 28:32]
  wire  fa_24_io_i0; // @[addsub.scala 28:32]
  wire  fa_24_io_i1; // @[addsub.scala 28:32]
  wire  fa_24_io_cin; // @[addsub.scala 28:32]
  wire  fa_24_io_sum; // @[addsub.scala 28:32]
  wire  fa_24_io_cout; // @[addsub.scala 28:32]
  wire  fa_25_io_i0; // @[addsub.scala 28:32]
  wire  fa_25_io_i1; // @[addsub.scala 28:32]
  wire  fa_25_io_cin; // @[addsub.scala 28:32]
  wire  fa_25_io_sum; // @[addsub.scala 28:32]
  wire  fa_25_io_cout; // @[addsub.scala 28:32]
  wire  fa_26_io_i0; // @[addsub.scala 28:32]
  wire  fa_26_io_i1; // @[addsub.scala 28:32]
  wire  fa_26_io_cin; // @[addsub.scala 28:32]
  wire  fa_26_io_sum; // @[addsub.scala 28:32]
  wire  fa_26_io_cout; // @[addsub.scala 28:32]
  wire  fa_27_io_i0; // @[addsub.scala 28:32]
  wire  fa_27_io_i1; // @[addsub.scala 28:32]
  wire  fa_27_io_cin; // @[addsub.scala 28:32]
  wire  fa_27_io_sum; // @[addsub.scala 28:32]
  wire  fa_27_io_cout; // @[addsub.scala 28:32]
  wire  fa_28_io_i0; // @[addsub.scala 28:32]
  wire  fa_28_io_i1; // @[addsub.scala 28:32]
  wire  fa_28_io_cin; // @[addsub.scala 28:32]
  wire  fa_28_io_sum; // @[addsub.scala 28:32]
  wire  fa_28_io_cout; // @[addsub.scala 28:32]
  wire  fa_29_io_i0; // @[addsub.scala 28:32]
  wire  fa_29_io_i1; // @[addsub.scala 28:32]
  wire  fa_29_io_cin; // @[addsub.scala 28:32]
  wire  fa_29_io_sum; // @[addsub.scala 28:32]
  wire  fa_29_io_cout; // @[addsub.scala 28:32]
  wire  fa_30_io_i0; // @[addsub.scala 28:32]
  wire  fa_30_io_i1; // @[addsub.scala 28:32]
  wire  fa_30_io_cin; // @[addsub.scala 28:32]
  wire  fa_30_io_sum; // @[addsub.scala 28:32]
  wire  fa_30_io_cout; // @[addsub.scala 28:32]
  wire  fa_31_io_i0; // @[addsub.scala 28:32]
  wire  fa_31_io_i1; // @[addsub.scala 28:32]
  wire  fa_31_io_cin; // @[addsub.scala 28:32]
  wire  fa_31_io_sum; // @[addsub.scala 28:32]
  wire  fa_31_io_cout; // @[addsub.scala 28:32]
  wire  fa_32_io_i0; // @[addsub.scala 28:32]
  wire  fa_32_io_i1; // @[addsub.scala 28:32]
  wire  fa_32_io_cin; // @[addsub.scala 28:32]
  wire  fa_32_io_sum; // @[addsub.scala 28:32]
  wire  fa_32_io_cout; // @[addsub.scala 28:32]
  wire  fa_33_io_i0; // @[addsub.scala 28:32]
  wire  fa_33_io_i1; // @[addsub.scala 28:32]
  wire  fa_33_io_cin; // @[addsub.scala 28:32]
  wire  fa_33_io_sum; // @[addsub.scala 28:32]
  wire  fa_33_io_cout; // @[addsub.scala 28:32]
  wire  fa_34_io_i0; // @[addsub.scala 28:32]
  wire  fa_34_io_i1; // @[addsub.scala 28:32]
  wire  fa_34_io_cin; // @[addsub.scala 28:32]
  wire  fa_34_io_sum; // @[addsub.scala 28:32]
  wire  fa_34_io_cout; // @[addsub.scala 28:32]
  wire  fa_35_io_i0; // @[addsub.scala 28:32]
  wire  fa_35_io_i1; // @[addsub.scala 28:32]
  wire  fa_35_io_cin; // @[addsub.scala 28:32]
  wire  fa_35_io_sum; // @[addsub.scala 28:32]
  wire  fa_35_io_cout; // @[addsub.scala 28:32]
  wire  fa_36_io_i0; // @[addsub.scala 28:32]
  wire  fa_36_io_i1; // @[addsub.scala 28:32]
  wire  fa_36_io_cin; // @[addsub.scala 28:32]
  wire  fa_36_io_sum; // @[addsub.scala 28:32]
  wire  fa_36_io_cout; // @[addsub.scala 28:32]
  wire  fa_37_io_i0; // @[addsub.scala 28:32]
  wire  fa_37_io_i1; // @[addsub.scala 28:32]
  wire  fa_37_io_cin; // @[addsub.scala 28:32]
  wire  fa_37_io_sum; // @[addsub.scala 28:32]
  wire  fa_37_io_cout; // @[addsub.scala 28:32]
  wire  fa_38_io_i0; // @[addsub.scala 28:32]
  wire  fa_38_io_i1; // @[addsub.scala 28:32]
  wire  fa_38_io_cin; // @[addsub.scala 28:32]
  wire  fa_38_io_sum; // @[addsub.scala 28:32]
  wire  fa_38_io_cout; // @[addsub.scala 28:32]
  wire  fa_39_io_i0; // @[addsub.scala 28:32]
  wire  fa_39_io_i1; // @[addsub.scala 28:32]
  wire  fa_39_io_cin; // @[addsub.scala 28:32]
  wire  fa_39_io_sum; // @[addsub.scala 28:32]
  wire  fa_39_io_cout; // @[addsub.scala 28:32]
  wire  fa_40_io_i0; // @[addsub.scala 28:32]
  wire  fa_40_io_i1; // @[addsub.scala 28:32]
  wire  fa_40_io_cin; // @[addsub.scala 28:32]
  wire  fa_40_io_sum; // @[addsub.scala 28:32]
  wire  fa_40_io_cout; // @[addsub.scala 28:32]
  wire  fa_41_io_i0; // @[addsub.scala 28:32]
  wire  fa_41_io_i1; // @[addsub.scala 28:32]
  wire  fa_41_io_cin; // @[addsub.scala 28:32]
  wire  fa_41_io_sum; // @[addsub.scala 28:32]
  wire  fa_41_io_cout; // @[addsub.scala 28:32]
  wire  fa_42_io_i0; // @[addsub.scala 28:32]
  wire  fa_42_io_i1; // @[addsub.scala 28:32]
  wire  fa_42_io_cin; // @[addsub.scala 28:32]
  wire  fa_42_io_sum; // @[addsub.scala 28:32]
  wire  fa_42_io_cout; // @[addsub.scala 28:32]
  wire  fa_43_io_i0; // @[addsub.scala 28:32]
  wire  fa_43_io_i1; // @[addsub.scala 28:32]
  wire  fa_43_io_cin; // @[addsub.scala 28:32]
  wire  fa_43_io_sum; // @[addsub.scala 28:32]
  wire  fa_43_io_cout; // @[addsub.scala 28:32]
  wire  fa_44_io_i0; // @[addsub.scala 28:32]
  wire  fa_44_io_i1; // @[addsub.scala 28:32]
  wire  fa_44_io_cin; // @[addsub.scala 28:32]
  wire  fa_44_io_sum; // @[addsub.scala 28:32]
  wire  fa_44_io_cout; // @[addsub.scala 28:32]
  wire  fa_45_io_i0; // @[addsub.scala 28:32]
  wire  fa_45_io_i1; // @[addsub.scala 28:32]
  wire  fa_45_io_cin; // @[addsub.scala 28:32]
  wire  fa_45_io_sum; // @[addsub.scala 28:32]
  wire  fa_45_io_cout; // @[addsub.scala 28:32]
  wire  fa_46_io_i0; // @[addsub.scala 28:32]
  wire  fa_46_io_i1; // @[addsub.scala 28:32]
  wire  fa_46_io_cin; // @[addsub.scala 28:32]
  wire  fa_46_io_sum; // @[addsub.scala 28:32]
  wire  fa_46_io_cout; // @[addsub.scala 28:32]
  wire  fa_47_io_i0; // @[addsub.scala 28:32]
  wire  fa_47_io_i1; // @[addsub.scala 28:32]
  wire  fa_47_io_cin; // @[addsub.scala 28:32]
  wire  fa_47_io_sum; // @[addsub.scala 28:32]
  wire  fa_47_io_cout; // @[addsub.scala 28:32]
  wire  fa_48_io_i0; // @[addsub.scala 28:32]
  wire  fa_48_io_i1; // @[addsub.scala 28:32]
  wire  fa_48_io_cin; // @[addsub.scala 28:32]
  wire  fa_48_io_sum; // @[addsub.scala 28:32]
  wire  fa_48_io_cout; // @[addsub.scala 28:32]
  wire  fa_49_io_i0; // @[addsub.scala 28:32]
  wire  fa_49_io_i1; // @[addsub.scala 28:32]
  wire  fa_49_io_cin; // @[addsub.scala 28:32]
  wire  fa_49_io_sum; // @[addsub.scala 28:32]
  wire  fa_49_io_cout; // @[addsub.scala 28:32]
  wire  fa_50_io_i0; // @[addsub.scala 28:32]
  wire  fa_50_io_i1; // @[addsub.scala 28:32]
  wire  fa_50_io_cin; // @[addsub.scala 28:32]
  wire  fa_50_io_sum; // @[addsub.scala 28:32]
  wire  fa_50_io_cout; // @[addsub.scala 28:32]
  wire  fa_51_io_i0; // @[addsub.scala 28:32]
  wire  fa_51_io_i1; // @[addsub.scala 28:32]
  wire  fa_51_io_cin; // @[addsub.scala 28:32]
  wire  fa_51_io_sum; // @[addsub.scala 28:32]
  wire  fa_51_io_cout; // @[addsub.scala 28:32]
  wire  fa_52_io_i0; // @[addsub.scala 28:32]
  wire  fa_52_io_i1; // @[addsub.scala 28:32]
  wire  fa_52_io_cin; // @[addsub.scala 28:32]
  wire  fa_52_io_sum; // @[addsub.scala 28:32]
  wire  fa_52_io_cout; // @[addsub.scala 28:32]
  wire  fa_53_io_i0; // @[addsub.scala 28:32]
  wire  fa_53_io_i1; // @[addsub.scala 28:32]
  wire  fa_53_io_cin; // @[addsub.scala 28:32]
  wire  fa_53_io_sum; // @[addsub.scala 28:32]
  wire  fa_53_io_cout; // @[addsub.scala 28:32]
  wire  fa_54_io_i0; // @[addsub.scala 28:32]
  wire  fa_54_io_i1; // @[addsub.scala 28:32]
  wire  fa_54_io_cin; // @[addsub.scala 28:32]
  wire  fa_54_io_sum; // @[addsub.scala 28:32]
  wire  fa_54_io_cout; // @[addsub.scala 28:32]
  wire  fa_55_io_i0; // @[addsub.scala 28:32]
  wire  fa_55_io_i1; // @[addsub.scala 28:32]
  wire  fa_55_io_cin; // @[addsub.scala 28:32]
  wire  fa_55_io_sum; // @[addsub.scala 28:32]
  wire  fa_55_io_cout; // @[addsub.scala 28:32]
  wire  fa_56_io_i0; // @[addsub.scala 28:32]
  wire  fa_56_io_i1; // @[addsub.scala 28:32]
  wire  fa_56_io_cin; // @[addsub.scala 28:32]
  wire  fa_56_io_sum; // @[addsub.scala 28:32]
  wire  fa_56_io_cout; // @[addsub.scala 28:32]
  wire  fa_57_io_i0; // @[addsub.scala 28:32]
  wire  fa_57_io_i1; // @[addsub.scala 28:32]
  wire  fa_57_io_cin; // @[addsub.scala 28:32]
  wire  fa_57_io_sum; // @[addsub.scala 28:32]
  wire  fa_57_io_cout; // @[addsub.scala 28:32]
  wire  fa_58_io_i0; // @[addsub.scala 28:32]
  wire  fa_58_io_i1; // @[addsub.scala 28:32]
  wire  fa_58_io_cin; // @[addsub.scala 28:32]
  wire  fa_58_io_sum; // @[addsub.scala 28:32]
  wire  fa_58_io_cout; // @[addsub.scala 28:32]
  wire  fa_59_io_i0; // @[addsub.scala 28:32]
  wire  fa_59_io_i1; // @[addsub.scala 28:32]
  wire  fa_59_io_cin; // @[addsub.scala 28:32]
  wire  fa_59_io_sum; // @[addsub.scala 28:32]
  wire  fa_59_io_cout; // @[addsub.scala 28:32]
  wire  fa_60_io_i0; // @[addsub.scala 28:32]
  wire  fa_60_io_i1; // @[addsub.scala 28:32]
  wire  fa_60_io_cin; // @[addsub.scala 28:32]
  wire  fa_60_io_sum; // @[addsub.scala 28:32]
  wire  fa_60_io_cout; // @[addsub.scala 28:32]
  wire  fa_61_io_i0; // @[addsub.scala 28:32]
  wire  fa_61_io_i1; // @[addsub.scala 28:32]
  wire  fa_61_io_cin; // @[addsub.scala 28:32]
  wire  fa_61_io_sum; // @[addsub.scala 28:32]
  wire  fa_61_io_cout; // @[addsub.scala 28:32]
  wire  fa_62_io_i0; // @[addsub.scala 28:32]
  wire  fa_62_io_i1; // @[addsub.scala 28:32]
  wire  fa_62_io_cin; // @[addsub.scala 28:32]
  wire  fa_62_io_sum; // @[addsub.scala 28:32]
  wire  fa_62_io_cout; // @[addsub.scala 28:32]
  wire  fa_63_io_i0; // @[addsub.scala 28:32]
  wire  fa_63_io_i1; // @[addsub.scala 28:32]
  wire  fa_63_io_cin; // @[addsub.scala 28:32]
  wire  fa_63_io_sum; // @[addsub.scala 28:32]
  wire  fa_63_io_cout; // @[addsub.scala 28:32]
  wire [7:0] lo_lo_lo = {fa_7_io_sum,fa_6_io_sum,fa_5_io_sum,fa_4_io_sum,fa_3_io_sum,fa_2_io_sum,fa_1_io_sum,fa_0_io_sum
    }; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {fa_15_io_sum,fa_14_io_sum,fa_13_io_sum,fa_12_io_sum,fa_11_io_sum,fa_10_io_sum,fa_9_io_sum,
    fa_8_io_sum,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {fa_23_io_sum,fa_22_io_sum,fa_21_io_sum,fa_20_io_sum,fa_19_io_sum,fa_18_io_sum,fa_17_io_sum,
    fa_16_io_sum}; // @[Cat.scala 30:58]
  wire [31:0] lo = {fa_31_io_sum,fa_30_io_sum,fa_29_io_sum,fa_28_io_sum,fa_27_io_sum,fa_26_io_sum,fa_25_io_sum,
    fa_24_io_sum,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {fa_39_io_sum,fa_38_io_sum,fa_37_io_sum,fa_36_io_sum,fa_35_io_sum,fa_34_io_sum,fa_33_io_sum,
    fa_32_io_sum}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {fa_47_io_sum,fa_46_io_sum,fa_45_io_sum,fa_44_io_sum,fa_43_io_sum,fa_42_io_sum,fa_41_io_sum,
    fa_40_io_sum,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {fa_55_io_sum,fa_54_io_sum,fa_53_io_sum,fa_52_io_sum,fa_51_io_sum,fa_50_io_sum,fa_49_io_sum,
    fa_48_io_sum}; // @[Cat.scala 30:58]
  wire [31:0] hi = {fa_63_io_sum,fa_62_io_sum,fa_61_io_sum,fa_60_io_sum,fa_59_io_sum,fa_58_io_sum,fa_57_io_sum,
    fa_56_io_sum,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  fullAdder fa_0 ( // @[addsub.scala 28:32]
    .io_i0(fa_0_io_i0),
    .io_i1(fa_0_io_i1),
    .io_cin(fa_0_io_cin),
    .io_sum(fa_0_io_sum),
    .io_cout(fa_0_io_cout)
  );
  fullAdder fa_1 ( // @[addsub.scala 28:32]
    .io_i0(fa_1_io_i0),
    .io_i1(fa_1_io_i1),
    .io_cin(fa_1_io_cin),
    .io_sum(fa_1_io_sum),
    .io_cout(fa_1_io_cout)
  );
  fullAdder fa_2 ( // @[addsub.scala 28:32]
    .io_i0(fa_2_io_i0),
    .io_i1(fa_2_io_i1),
    .io_cin(fa_2_io_cin),
    .io_sum(fa_2_io_sum),
    .io_cout(fa_2_io_cout)
  );
  fullAdder fa_3 ( // @[addsub.scala 28:32]
    .io_i0(fa_3_io_i0),
    .io_i1(fa_3_io_i1),
    .io_cin(fa_3_io_cin),
    .io_sum(fa_3_io_sum),
    .io_cout(fa_3_io_cout)
  );
  fullAdder fa_4 ( // @[addsub.scala 28:32]
    .io_i0(fa_4_io_i0),
    .io_i1(fa_4_io_i1),
    .io_cin(fa_4_io_cin),
    .io_sum(fa_4_io_sum),
    .io_cout(fa_4_io_cout)
  );
  fullAdder fa_5 ( // @[addsub.scala 28:32]
    .io_i0(fa_5_io_i0),
    .io_i1(fa_5_io_i1),
    .io_cin(fa_5_io_cin),
    .io_sum(fa_5_io_sum),
    .io_cout(fa_5_io_cout)
  );
  fullAdder fa_6 ( // @[addsub.scala 28:32]
    .io_i0(fa_6_io_i0),
    .io_i1(fa_6_io_i1),
    .io_cin(fa_6_io_cin),
    .io_sum(fa_6_io_sum),
    .io_cout(fa_6_io_cout)
  );
  fullAdder fa_7 ( // @[addsub.scala 28:32]
    .io_i0(fa_7_io_i0),
    .io_i1(fa_7_io_i1),
    .io_cin(fa_7_io_cin),
    .io_sum(fa_7_io_sum),
    .io_cout(fa_7_io_cout)
  );
  fullAdder fa_8 ( // @[addsub.scala 28:32]
    .io_i0(fa_8_io_i0),
    .io_i1(fa_8_io_i1),
    .io_cin(fa_8_io_cin),
    .io_sum(fa_8_io_sum),
    .io_cout(fa_8_io_cout)
  );
  fullAdder fa_9 ( // @[addsub.scala 28:32]
    .io_i0(fa_9_io_i0),
    .io_i1(fa_9_io_i1),
    .io_cin(fa_9_io_cin),
    .io_sum(fa_9_io_sum),
    .io_cout(fa_9_io_cout)
  );
  fullAdder fa_10 ( // @[addsub.scala 28:32]
    .io_i0(fa_10_io_i0),
    .io_i1(fa_10_io_i1),
    .io_cin(fa_10_io_cin),
    .io_sum(fa_10_io_sum),
    .io_cout(fa_10_io_cout)
  );
  fullAdder fa_11 ( // @[addsub.scala 28:32]
    .io_i0(fa_11_io_i0),
    .io_i1(fa_11_io_i1),
    .io_cin(fa_11_io_cin),
    .io_sum(fa_11_io_sum),
    .io_cout(fa_11_io_cout)
  );
  fullAdder fa_12 ( // @[addsub.scala 28:32]
    .io_i0(fa_12_io_i0),
    .io_i1(fa_12_io_i1),
    .io_cin(fa_12_io_cin),
    .io_sum(fa_12_io_sum),
    .io_cout(fa_12_io_cout)
  );
  fullAdder fa_13 ( // @[addsub.scala 28:32]
    .io_i0(fa_13_io_i0),
    .io_i1(fa_13_io_i1),
    .io_cin(fa_13_io_cin),
    .io_sum(fa_13_io_sum),
    .io_cout(fa_13_io_cout)
  );
  fullAdder fa_14 ( // @[addsub.scala 28:32]
    .io_i0(fa_14_io_i0),
    .io_i1(fa_14_io_i1),
    .io_cin(fa_14_io_cin),
    .io_sum(fa_14_io_sum),
    .io_cout(fa_14_io_cout)
  );
  fullAdder fa_15 ( // @[addsub.scala 28:32]
    .io_i0(fa_15_io_i0),
    .io_i1(fa_15_io_i1),
    .io_cin(fa_15_io_cin),
    .io_sum(fa_15_io_sum),
    .io_cout(fa_15_io_cout)
  );
  fullAdder fa_16 ( // @[addsub.scala 28:32]
    .io_i0(fa_16_io_i0),
    .io_i1(fa_16_io_i1),
    .io_cin(fa_16_io_cin),
    .io_sum(fa_16_io_sum),
    .io_cout(fa_16_io_cout)
  );
  fullAdder fa_17 ( // @[addsub.scala 28:32]
    .io_i0(fa_17_io_i0),
    .io_i1(fa_17_io_i1),
    .io_cin(fa_17_io_cin),
    .io_sum(fa_17_io_sum),
    .io_cout(fa_17_io_cout)
  );
  fullAdder fa_18 ( // @[addsub.scala 28:32]
    .io_i0(fa_18_io_i0),
    .io_i1(fa_18_io_i1),
    .io_cin(fa_18_io_cin),
    .io_sum(fa_18_io_sum),
    .io_cout(fa_18_io_cout)
  );
  fullAdder fa_19 ( // @[addsub.scala 28:32]
    .io_i0(fa_19_io_i0),
    .io_i1(fa_19_io_i1),
    .io_cin(fa_19_io_cin),
    .io_sum(fa_19_io_sum),
    .io_cout(fa_19_io_cout)
  );
  fullAdder fa_20 ( // @[addsub.scala 28:32]
    .io_i0(fa_20_io_i0),
    .io_i1(fa_20_io_i1),
    .io_cin(fa_20_io_cin),
    .io_sum(fa_20_io_sum),
    .io_cout(fa_20_io_cout)
  );
  fullAdder fa_21 ( // @[addsub.scala 28:32]
    .io_i0(fa_21_io_i0),
    .io_i1(fa_21_io_i1),
    .io_cin(fa_21_io_cin),
    .io_sum(fa_21_io_sum),
    .io_cout(fa_21_io_cout)
  );
  fullAdder fa_22 ( // @[addsub.scala 28:32]
    .io_i0(fa_22_io_i0),
    .io_i1(fa_22_io_i1),
    .io_cin(fa_22_io_cin),
    .io_sum(fa_22_io_sum),
    .io_cout(fa_22_io_cout)
  );
  fullAdder fa_23 ( // @[addsub.scala 28:32]
    .io_i0(fa_23_io_i0),
    .io_i1(fa_23_io_i1),
    .io_cin(fa_23_io_cin),
    .io_sum(fa_23_io_sum),
    .io_cout(fa_23_io_cout)
  );
  fullAdder fa_24 ( // @[addsub.scala 28:32]
    .io_i0(fa_24_io_i0),
    .io_i1(fa_24_io_i1),
    .io_cin(fa_24_io_cin),
    .io_sum(fa_24_io_sum),
    .io_cout(fa_24_io_cout)
  );
  fullAdder fa_25 ( // @[addsub.scala 28:32]
    .io_i0(fa_25_io_i0),
    .io_i1(fa_25_io_i1),
    .io_cin(fa_25_io_cin),
    .io_sum(fa_25_io_sum),
    .io_cout(fa_25_io_cout)
  );
  fullAdder fa_26 ( // @[addsub.scala 28:32]
    .io_i0(fa_26_io_i0),
    .io_i1(fa_26_io_i1),
    .io_cin(fa_26_io_cin),
    .io_sum(fa_26_io_sum),
    .io_cout(fa_26_io_cout)
  );
  fullAdder fa_27 ( // @[addsub.scala 28:32]
    .io_i0(fa_27_io_i0),
    .io_i1(fa_27_io_i1),
    .io_cin(fa_27_io_cin),
    .io_sum(fa_27_io_sum),
    .io_cout(fa_27_io_cout)
  );
  fullAdder fa_28 ( // @[addsub.scala 28:32]
    .io_i0(fa_28_io_i0),
    .io_i1(fa_28_io_i1),
    .io_cin(fa_28_io_cin),
    .io_sum(fa_28_io_sum),
    .io_cout(fa_28_io_cout)
  );
  fullAdder fa_29 ( // @[addsub.scala 28:32]
    .io_i0(fa_29_io_i0),
    .io_i1(fa_29_io_i1),
    .io_cin(fa_29_io_cin),
    .io_sum(fa_29_io_sum),
    .io_cout(fa_29_io_cout)
  );
  fullAdder fa_30 ( // @[addsub.scala 28:32]
    .io_i0(fa_30_io_i0),
    .io_i1(fa_30_io_i1),
    .io_cin(fa_30_io_cin),
    .io_sum(fa_30_io_sum),
    .io_cout(fa_30_io_cout)
  );
  fullAdder fa_31 ( // @[addsub.scala 28:32]
    .io_i0(fa_31_io_i0),
    .io_i1(fa_31_io_i1),
    .io_cin(fa_31_io_cin),
    .io_sum(fa_31_io_sum),
    .io_cout(fa_31_io_cout)
  );
  fullAdder fa_32 ( // @[addsub.scala 28:32]
    .io_i0(fa_32_io_i0),
    .io_i1(fa_32_io_i1),
    .io_cin(fa_32_io_cin),
    .io_sum(fa_32_io_sum),
    .io_cout(fa_32_io_cout)
  );
  fullAdder fa_33 ( // @[addsub.scala 28:32]
    .io_i0(fa_33_io_i0),
    .io_i1(fa_33_io_i1),
    .io_cin(fa_33_io_cin),
    .io_sum(fa_33_io_sum),
    .io_cout(fa_33_io_cout)
  );
  fullAdder fa_34 ( // @[addsub.scala 28:32]
    .io_i0(fa_34_io_i0),
    .io_i1(fa_34_io_i1),
    .io_cin(fa_34_io_cin),
    .io_sum(fa_34_io_sum),
    .io_cout(fa_34_io_cout)
  );
  fullAdder fa_35 ( // @[addsub.scala 28:32]
    .io_i0(fa_35_io_i0),
    .io_i1(fa_35_io_i1),
    .io_cin(fa_35_io_cin),
    .io_sum(fa_35_io_sum),
    .io_cout(fa_35_io_cout)
  );
  fullAdder fa_36 ( // @[addsub.scala 28:32]
    .io_i0(fa_36_io_i0),
    .io_i1(fa_36_io_i1),
    .io_cin(fa_36_io_cin),
    .io_sum(fa_36_io_sum),
    .io_cout(fa_36_io_cout)
  );
  fullAdder fa_37 ( // @[addsub.scala 28:32]
    .io_i0(fa_37_io_i0),
    .io_i1(fa_37_io_i1),
    .io_cin(fa_37_io_cin),
    .io_sum(fa_37_io_sum),
    .io_cout(fa_37_io_cout)
  );
  fullAdder fa_38 ( // @[addsub.scala 28:32]
    .io_i0(fa_38_io_i0),
    .io_i1(fa_38_io_i1),
    .io_cin(fa_38_io_cin),
    .io_sum(fa_38_io_sum),
    .io_cout(fa_38_io_cout)
  );
  fullAdder fa_39 ( // @[addsub.scala 28:32]
    .io_i0(fa_39_io_i0),
    .io_i1(fa_39_io_i1),
    .io_cin(fa_39_io_cin),
    .io_sum(fa_39_io_sum),
    .io_cout(fa_39_io_cout)
  );
  fullAdder fa_40 ( // @[addsub.scala 28:32]
    .io_i0(fa_40_io_i0),
    .io_i1(fa_40_io_i1),
    .io_cin(fa_40_io_cin),
    .io_sum(fa_40_io_sum),
    .io_cout(fa_40_io_cout)
  );
  fullAdder fa_41 ( // @[addsub.scala 28:32]
    .io_i0(fa_41_io_i0),
    .io_i1(fa_41_io_i1),
    .io_cin(fa_41_io_cin),
    .io_sum(fa_41_io_sum),
    .io_cout(fa_41_io_cout)
  );
  fullAdder fa_42 ( // @[addsub.scala 28:32]
    .io_i0(fa_42_io_i0),
    .io_i1(fa_42_io_i1),
    .io_cin(fa_42_io_cin),
    .io_sum(fa_42_io_sum),
    .io_cout(fa_42_io_cout)
  );
  fullAdder fa_43 ( // @[addsub.scala 28:32]
    .io_i0(fa_43_io_i0),
    .io_i1(fa_43_io_i1),
    .io_cin(fa_43_io_cin),
    .io_sum(fa_43_io_sum),
    .io_cout(fa_43_io_cout)
  );
  fullAdder fa_44 ( // @[addsub.scala 28:32]
    .io_i0(fa_44_io_i0),
    .io_i1(fa_44_io_i1),
    .io_cin(fa_44_io_cin),
    .io_sum(fa_44_io_sum),
    .io_cout(fa_44_io_cout)
  );
  fullAdder fa_45 ( // @[addsub.scala 28:32]
    .io_i0(fa_45_io_i0),
    .io_i1(fa_45_io_i1),
    .io_cin(fa_45_io_cin),
    .io_sum(fa_45_io_sum),
    .io_cout(fa_45_io_cout)
  );
  fullAdder fa_46 ( // @[addsub.scala 28:32]
    .io_i0(fa_46_io_i0),
    .io_i1(fa_46_io_i1),
    .io_cin(fa_46_io_cin),
    .io_sum(fa_46_io_sum),
    .io_cout(fa_46_io_cout)
  );
  fullAdder fa_47 ( // @[addsub.scala 28:32]
    .io_i0(fa_47_io_i0),
    .io_i1(fa_47_io_i1),
    .io_cin(fa_47_io_cin),
    .io_sum(fa_47_io_sum),
    .io_cout(fa_47_io_cout)
  );
  fullAdder fa_48 ( // @[addsub.scala 28:32]
    .io_i0(fa_48_io_i0),
    .io_i1(fa_48_io_i1),
    .io_cin(fa_48_io_cin),
    .io_sum(fa_48_io_sum),
    .io_cout(fa_48_io_cout)
  );
  fullAdder fa_49 ( // @[addsub.scala 28:32]
    .io_i0(fa_49_io_i0),
    .io_i1(fa_49_io_i1),
    .io_cin(fa_49_io_cin),
    .io_sum(fa_49_io_sum),
    .io_cout(fa_49_io_cout)
  );
  fullAdder fa_50 ( // @[addsub.scala 28:32]
    .io_i0(fa_50_io_i0),
    .io_i1(fa_50_io_i1),
    .io_cin(fa_50_io_cin),
    .io_sum(fa_50_io_sum),
    .io_cout(fa_50_io_cout)
  );
  fullAdder fa_51 ( // @[addsub.scala 28:32]
    .io_i0(fa_51_io_i0),
    .io_i1(fa_51_io_i1),
    .io_cin(fa_51_io_cin),
    .io_sum(fa_51_io_sum),
    .io_cout(fa_51_io_cout)
  );
  fullAdder fa_52 ( // @[addsub.scala 28:32]
    .io_i0(fa_52_io_i0),
    .io_i1(fa_52_io_i1),
    .io_cin(fa_52_io_cin),
    .io_sum(fa_52_io_sum),
    .io_cout(fa_52_io_cout)
  );
  fullAdder fa_53 ( // @[addsub.scala 28:32]
    .io_i0(fa_53_io_i0),
    .io_i1(fa_53_io_i1),
    .io_cin(fa_53_io_cin),
    .io_sum(fa_53_io_sum),
    .io_cout(fa_53_io_cout)
  );
  fullAdder fa_54 ( // @[addsub.scala 28:32]
    .io_i0(fa_54_io_i0),
    .io_i1(fa_54_io_i1),
    .io_cin(fa_54_io_cin),
    .io_sum(fa_54_io_sum),
    .io_cout(fa_54_io_cout)
  );
  fullAdder fa_55 ( // @[addsub.scala 28:32]
    .io_i0(fa_55_io_i0),
    .io_i1(fa_55_io_i1),
    .io_cin(fa_55_io_cin),
    .io_sum(fa_55_io_sum),
    .io_cout(fa_55_io_cout)
  );
  fullAdder fa_56 ( // @[addsub.scala 28:32]
    .io_i0(fa_56_io_i0),
    .io_i1(fa_56_io_i1),
    .io_cin(fa_56_io_cin),
    .io_sum(fa_56_io_sum),
    .io_cout(fa_56_io_cout)
  );
  fullAdder fa_57 ( // @[addsub.scala 28:32]
    .io_i0(fa_57_io_i0),
    .io_i1(fa_57_io_i1),
    .io_cin(fa_57_io_cin),
    .io_sum(fa_57_io_sum),
    .io_cout(fa_57_io_cout)
  );
  fullAdder fa_58 ( // @[addsub.scala 28:32]
    .io_i0(fa_58_io_i0),
    .io_i1(fa_58_io_i1),
    .io_cin(fa_58_io_cin),
    .io_sum(fa_58_io_sum),
    .io_cout(fa_58_io_cout)
  );
  fullAdder fa_59 ( // @[addsub.scala 28:32]
    .io_i0(fa_59_io_i0),
    .io_i1(fa_59_io_i1),
    .io_cin(fa_59_io_cin),
    .io_sum(fa_59_io_sum),
    .io_cout(fa_59_io_cout)
  );
  fullAdder fa_60 ( // @[addsub.scala 28:32]
    .io_i0(fa_60_io_i0),
    .io_i1(fa_60_io_i1),
    .io_cin(fa_60_io_cin),
    .io_sum(fa_60_io_sum),
    .io_cout(fa_60_io_cout)
  );
  fullAdder fa_61 ( // @[addsub.scala 28:32]
    .io_i0(fa_61_io_i0),
    .io_i1(fa_61_io_i1),
    .io_cin(fa_61_io_cin),
    .io_sum(fa_61_io_sum),
    .io_cout(fa_61_io_cout)
  );
  fullAdder fa_62 ( // @[addsub.scala 28:32]
    .io_i0(fa_62_io_i0),
    .io_i1(fa_62_io_i1),
    .io_cin(fa_62_io_cin),
    .io_sum(fa_62_io_sum),
    .io_cout(fa_62_io_cout)
  );
  fullAdder fa_63 ( // @[addsub.scala 28:32]
    .io_i0(fa_63_io_i0),
    .io_i1(fa_63_io_i1),
    .io_cin(fa_63_io_cin),
    .io_sum(fa_63_io_sum),
    .io_cout(fa_63_io_cout)
  );
  assign io_sum = {hi,lo}; // @[Cat.scala 30:58]
  assign fa_0_io_i0 = io_i0[0]; // @[addsub.scala 31:25]
  assign fa_0_io_i1 = io_onesComp_ip[0]; // @[addsub.scala 32:34]
  assign fa_0_io_cin = 1'h1; // @[addsub.scala 33:18]
  assign fa_1_io_i0 = io_i0[1]; // @[addsub.scala 37:29]
  assign fa_1_io_i1 = io_onesComp_ip[1]; // @[addsub.scala 38:38]
  assign fa_1_io_cin = fa_0_io_cout; // @[addsub.scala 39:22]
  assign fa_2_io_i0 = io_i0[2]; // @[addsub.scala 37:29]
  assign fa_2_io_i1 = io_onesComp_ip[2]; // @[addsub.scala 38:38]
  assign fa_2_io_cin = fa_1_io_cout; // @[addsub.scala 39:22]
  assign fa_3_io_i0 = io_i0[3]; // @[addsub.scala 37:29]
  assign fa_3_io_i1 = io_onesComp_ip[3]; // @[addsub.scala 38:38]
  assign fa_3_io_cin = fa_2_io_cout; // @[addsub.scala 39:22]
  assign fa_4_io_i0 = io_i0[4]; // @[addsub.scala 37:29]
  assign fa_4_io_i1 = io_onesComp_ip[4]; // @[addsub.scala 38:38]
  assign fa_4_io_cin = fa_3_io_cout; // @[addsub.scala 39:22]
  assign fa_5_io_i0 = io_i0[5]; // @[addsub.scala 37:29]
  assign fa_5_io_i1 = io_onesComp_ip[5]; // @[addsub.scala 38:38]
  assign fa_5_io_cin = fa_4_io_cout; // @[addsub.scala 39:22]
  assign fa_6_io_i0 = io_i0[6]; // @[addsub.scala 37:29]
  assign fa_6_io_i1 = io_onesComp_ip[6]; // @[addsub.scala 38:38]
  assign fa_6_io_cin = fa_5_io_cout; // @[addsub.scala 39:22]
  assign fa_7_io_i0 = io_i0[7]; // @[addsub.scala 37:29]
  assign fa_7_io_i1 = io_onesComp_ip[7]; // @[addsub.scala 38:38]
  assign fa_7_io_cin = fa_6_io_cout; // @[addsub.scala 39:22]
  assign fa_8_io_i0 = io_i0[8]; // @[addsub.scala 37:29]
  assign fa_8_io_i1 = io_onesComp_ip[8]; // @[addsub.scala 38:38]
  assign fa_8_io_cin = fa_7_io_cout; // @[addsub.scala 39:22]
  assign fa_9_io_i0 = io_i0[9]; // @[addsub.scala 37:29]
  assign fa_9_io_i1 = io_onesComp_ip[9]; // @[addsub.scala 38:38]
  assign fa_9_io_cin = fa_8_io_cout; // @[addsub.scala 39:22]
  assign fa_10_io_i0 = io_i0[10]; // @[addsub.scala 37:29]
  assign fa_10_io_i1 = io_onesComp_ip[10]; // @[addsub.scala 38:38]
  assign fa_10_io_cin = fa_9_io_cout; // @[addsub.scala 39:22]
  assign fa_11_io_i0 = io_i0[11]; // @[addsub.scala 37:29]
  assign fa_11_io_i1 = io_onesComp_ip[11]; // @[addsub.scala 38:38]
  assign fa_11_io_cin = fa_10_io_cout; // @[addsub.scala 39:22]
  assign fa_12_io_i0 = io_i0[12]; // @[addsub.scala 37:29]
  assign fa_12_io_i1 = io_onesComp_ip[12]; // @[addsub.scala 38:38]
  assign fa_12_io_cin = fa_11_io_cout; // @[addsub.scala 39:22]
  assign fa_13_io_i0 = io_i0[13]; // @[addsub.scala 37:29]
  assign fa_13_io_i1 = io_onesComp_ip[13]; // @[addsub.scala 38:38]
  assign fa_13_io_cin = fa_12_io_cout; // @[addsub.scala 39:22]
  assign fa_14_io_i0 = io_i0[14]; // @[addsub.scala 37:29]
  assign fa_14_io_i1 = io_onesComp_ip[14]; // @[addsub.scala 38:38]
  assign fa_14_io_cin = fa_13_io_cout; // @[addsub.scala 39:22]
  assign fa_15_io_i0 = io_i0[15]; // @[addsub.scala 37:29]
  assign fa_15_io_i1 = io_onesComp_ip[15]; // @[addsub.scala 38:38]
  assign fa_15_io_cin = fa_14_io_cout; // @[addsub.scala 39:22]
  assign fa_16_io_i0 = io_i0[16]; // @[addsub.scala 37:29]
  assign fa_16_io_i1 = io_onesComp_ip[16]; // @[addsub.scala 38:38]
  assign fa_16_io_cin = fa_15_io_cout; // @[addsub.scala 39:22]
  assign fa_17_io_i0 = io_i0[17]; // @[addsub.scala 37:29]
  assign fa_17_io_i1 = io_onesComp_ip[17]; // @[addsub.scala 38:38]
  assign fa_17_io_cin = fa_16_io_cout; // @[addsub.scala 39:22]
  assign fa_18_io_i0 = io_i0[18]; // @[addsub.scala 37:29]
  assign fa_18_io_i1 = io_onesComp_ip[18]; // @[addsub.scala 38:38]
  assign fa_18_io_cin = fa_17_io_cout; // @[addsub.scala 39:22]
  assign fa_19_io_i0 = io_i0[19]; // @[addsub.scala 37:29]
  assign fa_19_io_i1 = io_onesComp_ip[19]; // @[addsub.scala 38:38]
  assign fa_19_io_cin = fa_18_io_cout; // @[addsub.scala 39:22]
  assign fa_20_io_i0 = io_i0[20]; // @[addsub.scala 37:29]
  assign fa_20_io_i1 = io_onesComp_ip[20]; // @[addsub.scala 38:38]
  assign fa_20_io_cin = fa_19_io_cout; // @[addsub.scala 39:22]
  assign fa_21_io_i0 = io_i0[21]; // @[addsub.scala 37:29]
  assign fa_21_io_i1 = io_onesComp_ip[21]; // @[addsub.scala 38:38]
  assign fa_21_io_cin = fa_20_io_cout; // @[addsub.scala 39:22]
  assign fa_22_io_i0 = io_i0[22]; // @[addsub.scala 37:29]
  assign fa_22_io_i1 = io_onesComp_ip[22]; // @[addsub.scala 38:38]
  assign fa_22_io_cin = fa_21_io_cout; // @[addsub.scala 39:22]
  assign fa_23_io_i0 = io_i0[23]; // @[addsub.scala 37:29]
  assign fa_23_io_i1 = io_onesComp_ip[23]; // @[addsub.scala 38:38]
  assign fa_23_io_cin = fa_22_io_cout; // @[addsub.scala 39:22]
  assign fa_24_io_i0 = io_i0[24]; // @[addsub.scala 37:29]
  assign fa_24_io_i1 = io_onesComp_ip[24]; // @[addsub.scala 38:38]
  assign fa_24_io_cin = fa_23_io_cout; // @[addsub.scala 39:22]
  assign fa_25_io_i0 = io_i0[25]; // @[addsub.scala 37:29]
  assign fa_25_io_i1 = io_onesComp_ip[25]; // @[addsub.scala 38:38]
  assign fa_25_io_cin = fa_24_io_cout; // @[addsub.scala 39:22]
  assign fa_26_io_i0 = io_i0[26]; // @[addsub.scala 37:29]
  assign fa_26_io_i1 = io_onesComp_ip[26]; // @[addsub.scala 38:38]
  assign fa_26_io_cin = fa_25_io_cout; // @[addsub.scala 39:22]
  assign fa_27_io_i0 = io_i0[27]; // @[addsub.scala 37:29]
  assign fa_27_io_i1 = io_onesComp_ip[27]; // @[addsub.scala 38:38]
  assign fa_27_io_cin = fa_26_io_cout; // @[addsub.scala 39:22]
  assign fa_28_io_i0 = io_i0[28]; // @[addsub.scala 37:29]
  assign fa_28_io_i1 = io_onesComp_ip[28]; // @[addsub.scala 38:38]
  assign fa_28_io_cin = fa_27_io_cout; // @[addsub.scala 39:22]
  assign fa_29_io_i0 = io_i0[29]; // @[addsub.scala 37:29]
  assign fa_29_io_i1 = io_onesComp_ip[29]; // @[addsub.scala 38:38]
  assign fa_29_io_cin = fa_28_io_cout; // @[addsub.scala 39:22]
  assign fa_30_io_i0 = io_i0[30]; // @[addsub.scala 37:29]
  assign fa_30_io_i1 = io_onesComp_ip[30]; // @[addsub.scala 38:38]
  assign fa_30_io_cin = fa_29_io_cout; // @[addsub.scala 39:22]
  assign fa_31_io_i0 = io_i0[31]; // @[addsub.scala 37:29]
  assign fa_31_io_i1 = io_onesComp_ip[31]; // @[addsub.scala 38:38]
  assign fa_31_io_cin = fa_30_io_cout; // @[addsub.scala 39:22]
  assign fa_32_io_i0 = io_i0[32]; // @[addsub.scala 37:29]
  assign fa_32_io_i1 = io_onesComp_ip[32]; // @[addsub.scala 38:38]
  assign fa_32_io_cin = fa_31_io_cout; // @[addsub.scala 39:22]
  assign fa_33_io_i0 = io_i0[33]; // @[addsub.scala 37:29]
  assign fa_33_io_i1 = io_onesComp_ip[33]; // @[addsub.scala 38:38]
  assign fa_33_io_cin = fa_32_io_cout; // @[addsub.scala 39:22]
  assign fa_34_io_i0 = io_i0[34]; // @[addsub.scala 37:29]
  assign fa_34_io_i1 = io_onesComp_ip[34]; // @[addsub.scala 38:38]
  assign fa_34_io_cin = fa_33_io_cout; // @[addsub.scala 39:22]
  assign fa_35_io_i0 = io_i0[35]; // @[addsub.scala 37:29]
  assign fa_35_io_i1 = io_onesComp_ip[35]; // @[addsub.scala 38:38]
  assign fa_35_io_cin = fa_34_io_cout; // @[addsub.scala 39:22]
  assign fa_36_io_i0 = io_i0[36]; // @[addsub.scala 37:29]
  assign fa_36_io_i1 = io_onesComp_ip[36]; // @[addsub.scala 38:38]
  assign fa_36_io_cin = fa_35_io_cout; // @[addsub.scala 39:22]
  assign fa_37_io_i0 = io_i0[37]; // @[addsub.scala 37:29]
  assign fa_37_io_i1 = io_onesComp_ip[37]; // @[addsub.scala 38:38]
  assign fa_37_io_cin = fa_36_io_cout; // @[addsub.scala 39:22]
  assign fa_38_io_i0 = io_i0[38]; // @[addsub.scala 37:29]
  assign fa_38_io_i1 = io_onesComp_ip[38]; // @[addsub.scala 38:38]
  assign fa_38_io_cin = fa_37_io_cout; // @[addsub.scala 39:22]
  assign fa_39_io_i0 = io_i0[39]; // @[addsub.scala 37:29]
  assign fa_39_io_i1 = io_onesComp_ip[39]; // @[addsub.scala 38:38]
  assign fa_39_io_cin = fa_38_io_cout; // @[addsub.scala 39:22]
  assign fa_40_io_i0 = io_i0[40]; // @[addsub.scala 37:29]
  assign fa_40_io_i1 = io_onesComp_ip[40]; // @[addsub.scala 38:38]
  assign fa_40_io_cin = fa_39_io_cout; // @[addsub.scala 39:22]
  assign fa_41_io_i0 = io_i0[41]; // @[addsub.scala 37:29]
  assign fa_41_io_i1 = io_onesComp_ip[41]; // @[addsub.scala 38:38]
  assign fa_41_io_cin = fa_40_io_cout; // @[addsub.scala 39:22]
  assign fa_42_io_i0 = io_i0[42]; // @[addsub.scala 37:29]
  assign fa_42_io_i1 = io_onesComp_ip[42]; // @[addsub.scala 38:38]
  assign fa_42_io_cin = fa_41_io_cout; // @[addsub.scala 39:22]
  assign fa_43_io_i0 = io_i0[43]; // @[addsub.scala 37:29]
  assign fa_43_io_i1 = io_onesComp_ip[43]; // @[addsub.scala 38:38]
  assign fa_43_io_cin = fa_42_io_cout; // @[addsub.scala 39:22]
  assign fa_44_io_i0 = io_i0[44]; // @[addsub.scala 37:29]
  assign fa_44_io_i1 = io_onesComp_ip[44]; // @[addsub.scala 38:38]
  assign fa_44_io_cin = fa_43_io_cout; // @[addsub.scala 39:22]
  assign fa_45_io_i0 = io_i0[45]; // @[addsub.scala 37:29]
  assign fa_45_io_i1 = io_onesComp_ip[45]; // @[addsub.scala 38:38]
  assign fa_45_io_cin = fa_44_io_cout; // @[addsub.scala 39:22]
  assign fa_46_io_i0 = io_i0[46]; // @[addsub.scala 37:29]
  assign fa_46_io_i1 = io_onesComp_ip[46]; // @[addsub.scala 38:38]
  assign fa_46_io_cin = fa_45_io_cout; // @[addsub.scala 39:22]
  assign fa_47_io_i0 = io_i0[47]; // @[addsub.scala 37:29]
  assign fa_47_io_i1 = io_onesComp_ip[47]; // @[addsub.scala 38:38]
  assign fa_47_io_cin = fa_46_io_cout; // @[addsub.scala 39:22]
  assign fa_48_io_i0 = io_i0[48]; // @[addsub.scala 37:29]
  assign fa_48_io_i1 = io_onesComp_ip[48]; // @[addsub.scala 38:38]
  assign fa_48_io_cin = fa_47_io_cout; // @[addsub.scala 39:22]
  assign fa_49_io_i0 = io_i0[49]; // @[addsub.scala 37:29]
  assign fa_49_io_i1 = io_onesComp_ip[49]; // @[addsub.scala 38:38]
  assign fa_49_io_cin = fa_48_io_cout; // @[addsub.scala 39:22]
  assign fa_50_io_i0 = io_i0[50]; // @[addsub.scala 37:29]
  assign fa_50_io_i1 = io_onesComp_ip[50]; // @[addsub.scala 38:38]
  assign fa_50_io_cin = fa_49_io_cout; // @[addsub.scala 39:22]
  assign fa_51_io_i0 = io_i0[51]; // @[addsub.scala 37:29]
  assign fa_51_io_i1 = io_onesComp_ip[51]; // @[addsub.scala 38:38]
  assign fa_51_io_cin = fa_50_io_cout; // @[addsub.scala 39:22]
  assign fa_52_io_i0 = io_i0[52]; // @[addsub.scala 37:29]
  assign fa_52_io_i1 = io_onesComp_ip[52]; // @[addsub.scala 38:38]
  assign fa_52_io_cin = fa_51_io_cout; // @[addsub.scala 39:22]
  assign fa_53_io_i0 = io_i0[53]; // @[addsub.scala 37:29]
  assign fa_53_io_i1 = io_onesComp_ip[53]; // @[addsub.scala 38:38]
  assign fa_53_io_cin = fa_52_io_cout; // @[addsub.scala 39:22]
  assign fa_54_io_i0 = io_i0[54]; // @[addsub.scala 37:29]
  assign fa_54_io_i1 = io_onesComp_ip[54]; // @[addsub.scala 38:38]
  assign fa_54_io_cin = fa_53_io_cout; // @[addsub.scala 39:22]
  assign fa_55_io_i0 = io_i0[55]; // @[addsub.scala 37:29]
  assign fa_55_io_i1 = io_onesComp_ip[55]; // @[addsub.scala 38:38]
  assign fa_55_io_cin = fa_54_io_cout; // @[addsub.scala 39:22]
  assign fa_56_io_i0 = io_i0[56]; // @[addsub.scala 37:29]
  assign fa_56_io_i1 = io_onesComp_ip[56]; // @[addsub.scala 38:38]
  assign fa_56_io_cin = fa_55_io_cout; // @[addsub.scala 39:22]
  assign fa_57_io_i0 = io_i0[57]; // @[addsub.scala 37:29]
  assign fa_57_io_i1 = io_onesComp_ip[57]; // @[addsub.scala 38:38]
  assign fa_57_io_cin = fa_56_io_cout; // @[addsub.scala 39:22]
  assign fa_58_io_i0 = io_i0[58]; // @[addsub.scala 37:29]
  assign fa_58_io_i1 = io_onesComp_ip[58]; // @[addsub.scala 38:38]
  assign fa_58_io_cin = fa_57_io_cout; // @[addsub.scala 39:22]
  assign fa_59_io_i0 = io_i0[59]; // @[addsub.scala 37:29]
  assign fa_59_io_i1 = io_onesComp_ip[59]; // @[addsub.scala 38:38]
  assign fa_59_io_cin = fa_58_io_cout; // @[addsub.scala 39:22]
  assign fa_60_io_i0 = io_i0[60]; // @[addsub.scala 37:29]
  assign fa_60_io_i1 = io_onesComp_ip[60]; // @[addsub.scala 38:38]
  assign fa_60_io_cin = fa_59_io_cout; // @[addsub.scala 39:22]
  assign fa_61_io_i0 = io_i0[61]; // @[addsub.scala 37:29]
  assign fa_61_io_i1 = io_onesComp_ip[61]; // @[addsub.scala 38:38]
  assign fa_61_io_cin = fa_60_io_cout; // @[addsub.scala 39:22]
  assign fa_62_io_i0 = io_i0[62]; // @[addsub.scala 37:29]
  assign fa_62_io_i1 = io_onesComp_ip[62]; // @[addsub.scala 38:38]
  assign fa_62_io_cin = fa_61_io_cout; // @[addsub.scala 39:22]
  assign fa_63_io_i0 = io_i0[63]; // @[addsub.scala 37:29]
  assign fa_63_io_i1 = io_onesComp_ip[63]; // @[addsub.scala 38:38]
  assign fa_63_io_cin = fa_62_io_cout; // @[addsub.scala 39:22]
endmodule
module booth_div_substep(
  input  [63:0] io_acc,
  input  [63:0] io_Q,
  input  [63:0] io_divisor,
  output [63:0] io_next_acc,
  output [63:0] io_next_Q
);
  wire [63:0] g1_io_i1; // @[booth_div_substep.scala 13:20]
  wire [63:0] g1_io_onesComp; // @[booth_div_substep.scala 13:20]
  wire [63:0] as1_io_onesComp_ip; // @[booth_div_substep.scala 32:21]
  wire [63:0] as1_io_i0; // @[booth_div_substep.scala 32:21]
  wire [63:0] as1_io_sum; // @[booth_div_substep.scala 32:21]
  wire [64:0] shiftedA = {io_acc, 1'h0}; // @[booth_div_substep.scala 28:24]
  wire [64:0] shiftedQ = {io_Q, 1'h0}; // @[booth_div_substep.scala 30:22]
  wire [62:0] hi = shiftedA[63:1]; // @[booth_div_substep.scala 38:30]
  wire [64:0] shiftedA_LSB = {{64'd0}, io_Q[63]}; // @[booth_div_substep.scala 24:28 booth_div_substep.scala 29:18]
  wire [127:0] _T_3 = {hi,shiftedA_LSB}; // @[Cat.scala 30:58]
  wire [63:0] sub_temp = as1_io_sum; // @[booth_div_substep.scala 34:24 booth_div_substep.scala 39:14]
  wire  _GEN_0 = sub_temp[63] ? 1'h0 : 1'h1; // @[booth_div_substep.scala 42:33 booth_div_substep.scala 43:22 booth_div_substep.scala 46:22]
  wire [127:0] _GEN_1 = sub_temp[63] ? _T_3 : {{64'd0}, sub_temp}; // @[booth_div_substep.scala 42:33 booth_div_substep.scala 44:22 booth_div_substep.scala 47:22]
  wire [62:0] hi_2 = shiftedQ[63:1]; // @[booth_div_substep.scala 51:32]
  wire [64:0] shiftedQ_LSB = {{64'd0}, _GEN_0}; // @[booth_div_substep.scala 25:28]
  wire [127:0] _T_7 = {hi_2,shiftedQ_LSB}; // @[Cat.scala 30:58]
  wire [64:0] Aout = _GEN_1[64:0]; // @[booth_div_substep.scala 26:20]
  getOnesComplement g1 ( // @[booth_div_substep.scala 13:20]
    .io_i1(g1_io_i1),
    .io_onesComp(g1_io_onesComp)
  );
  addsub as1 ( // @[booth_div_substep.scala 32:21]
    .io_onesComp_ip(as1_io_onesComp_ip),
    .io_i0(as1_io_i0),
    .io_sum(as1_io_sum)
  );
  assign io_next_acc = Aout[63:0]; // @[booth_div_substep.scala 50:17]
  assign io_next_Q = _T_7[63:0]; // @[booth_div_substep.scala 51:17]
  assign g1_io_i1 = io_divisor; // @[booth_div_substep.scala 18:14]
  assign as1_io_onesComp_ip = g1_io_onesComp; // @[booth_div_substep.scala 15:22 booth_div_substep.scala 19:12]
  assign as1_io_i0 = _T_3[63:0]; // @[booth_div_substep.scala 38:15]
endmodule
module booth_divider(
  input         clock,
  input         reset,
  input         io_signed,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  output [63:0] io_quotient,
  output [63:0] io_remainder
);
  wire [63:0] bds_0_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_0_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_0_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_0_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_0_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_1_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_1_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_1_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_1_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_1_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_2_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_2_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_2_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_2_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_2_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_3_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_3_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_3_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_3_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_3_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_4_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_4_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_4_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_4_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_4_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_5_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_5_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_5_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_5_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_5_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_6_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_6_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_6_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_6_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_6_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_7_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_7_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_7_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_7_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_7_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_8_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_8_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_8_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_8_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_8_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_9_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_9_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_9_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_9_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_9_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_10_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_10_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_10_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_10_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_10_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_11_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_11_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_11_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_11_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_11_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_12_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_12_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_12_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_12_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_12_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_13_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_13_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_13_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_13_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_13_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_14_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_14_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_14_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_14_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_14_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_15_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_15_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_15_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_15_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_15_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_16_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_16_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_16_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_16_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_16_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_17_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_17_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_17_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_17_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_17_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_18_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_18_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_18_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_18_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_18_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_19_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_19_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_19_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_19_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_19_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_20_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_20_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_20_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_20_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_20_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_21_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_21_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_21_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_21_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_21_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_22_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_22_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_22_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_22_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_22_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_23_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_23_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_23_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_23_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_23_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_24_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_24_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_24_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_24_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_24_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_25_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_25_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_25_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_25_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_25_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_26_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_26_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_26_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_26_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_26_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_27_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_27_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_27_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_27_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_27_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_28_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_28_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_28_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_28_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_28_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_29_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_29_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_29_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_29_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_29_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_30_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_30_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_30_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_30_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_30_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_31_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_31_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_31_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_31_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_31_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_32_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_32_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_32_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_32_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_32_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_33_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_33_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_33_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_33_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_33_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_34_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_34_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_34_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_34_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_34_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_35_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_35_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_35_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_35_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_35_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_36_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_36_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_36_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_36_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_36_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_37_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_37_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_37_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_37_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_37_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_38_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_38_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_38_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_38_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_38_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_39_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_39_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_39_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_39_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_39_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_40_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_40_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_40_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_40_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_40_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_41_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_41_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_41_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_41_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_41_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_42_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_42_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_42_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_42_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_42_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_43_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_43_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_43_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_43_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_43_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_44_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_44_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_44_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_44_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_44_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_45_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_45_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_45_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_45_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_45_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_46_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_46_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_46_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_46_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_46_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_47_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_47_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_47_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_47_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_47_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_48_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_48_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_48_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_48_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_48_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_49_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_49_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_49_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_49_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_49_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_50_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_50_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_50_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_50_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_50_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_51_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_51_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_51_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_51_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_51_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_52_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_52_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_52_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_52_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_52_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_53_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_53_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_53_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_53_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_53_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_54_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_54_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_54_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_54_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_54_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_55_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_55_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_55_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_55_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_55_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_56_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_56_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_56_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_56_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_56_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_57_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_57_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_57_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_57_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_57_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_58_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_58_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_58_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_58_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_58_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_59_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_59_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_59_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_59_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_59_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_60_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_60_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_60_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_60_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_60_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_61_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_61_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_61_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_61_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_61_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_62_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_62_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_62_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_62_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_62_io_next_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_63_io_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_63_io_Q; // @[booth_divider.scala 51:33]
  wire [63:0] bds_63_io_divisor; // @[booth_divider.scala 51:33]
  wire [63:0] bds_63_io_next_acc; // @[booth_divider.scala 51:33]
  wire [63:0] bds_63_io_next_Q; // @[booth_divider.scala 51:33]
  wire  neg_quotient = (io_dividend[63] ^ io_divisor[63]) & io_signed; // @[booth_divider.scala 18:58]
  wire [63:0] _T_6 = ~io_dividend; // @[booth_divider.scala 24:22]
  wire [63:0] dividend_comp = _T_6 + 64'h1; // @[booth_divider.scala 24:42]
  wire [63:0] _T_10 = ~io_divisor; // @[booth_divider.scala 25:22]
  wire [63:0] divisor_comp = _T_10 + 64'h1; // @[booth_divider.scala 25:41]
  wire  _T_16 = io_signed & io_dividend[63]; // @[booth_divider.scala 29:29]
  wire [63:0] quotientTemp = bds_63_io_next_Q; // @[booth_divider.scala 45:29 booth_divider.scala 64:29]
  wire [63:0] _T_24 = ~quotientTemp; // @[booth_divider.scala 69:47]
  wire [63:0] _T_26 = _T_24 + 64'h1; // @[booth_divider.scala 69:61]
  wire [63:0] remainderTemp = bds_63_io_next_acc; // @[booth_divider.scala 46:29 booth_divider.scala 65:29]
  wire [63:0] _T_33 = ~remainderTemp; // @[booth_divider.scala 70:74]
  wire [63:0] _T_35 = _T_33 + 64'h1; // @[booth_divider.scala 70:89]
  booth_div_substep bds_0 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_0_io_acc),
    .io_Q(bds_0_io_Q),
    .io_divisor(bds_0_io_divisor),
    .io_next_acc(bds_0_io_next_acc),
    .io_next_Q(bds_0_io_next_Q)
  );
  booth_div_substep bds_1 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_1_io_acc),
    .io_Q(bds_1_io_Q),
    .io_divisor(bds_1_io_divisor),
    .io_next_acc(bds_1_io_next_acc),
    .io_next_Q(bds_1_io_next_Q)
  );
  booth_div_substep bds_2 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_2_io_acc),
    .io_Q(bds_2_io_Q),
    .io_divisor(bds_2_io_divisor),
    .io_next_acc(bds_2_io_next_acc),
    .io_next_Q(bds_2_io_next_Q)
  );
  booth_div_substep bds_3 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_3_io_acc),
    .io_Q(bds_3_io_Q),
    .io_divisor(bds_3_io_divisor),
    .io_next_acc(bds_3_io_next_acc),
    .io_next_Q(bds_3_io_next_Q)
  );
  booth_div_substep bds_4 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_4_io_acc),
    .io_Q(bds_4_io_Q),
    .io_divisor(bds_4_io_divisor),
    .io_next_acc(bds_4_io_next_acc),
    .io_next_Q(bds_4_io_next_Q)
  );
  booth_div_substep bds_5 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_5_io_acc),
    .io_Q(bds_5_io_Q),
    .io_divisor(bds_5_io_divisor),
    .io_next_acc(bds_5_io_next_acc),
    .io_next_Q(bds_5_io_next_Q)
  );
  booth_div_substep bds_6 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_6_io_acc),
    .io_Q(bds_6_io_Q),
    .io_divisor(bds_6_io_divisor),
    .io_next_acc(bds_6_io_next_acc),
    .io_next_Q(bds_6_io_next_Q)
  );
  booth_div_substep bds_7 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_7_io_acc),
    .io_Q(bds_7_io_Q),
    .io_divisor(bds_7_io_divisor),
    .io_next_acc(bds_7_io_next_acc),
    .io_next_Q(bds_7_io_next_Q)
  );
  booth_div_substep bds_8 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_8_io_acc),
    .io_Q(bds_8_io_Q),
    .io_divisor(bds_8_io_divisor),
    .io_next_acc(bds_8_io_next_acc),
    .io_next_Q(bds_8_io_next_Q)
  );
  booth_div_substep bds_9 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_9_io_acc),
    .io_Q(bds_9_io_Q),
    .io_divisor(bds_9_io_divisor),
    .io_next_acc(bds_9_io_next_acc),
    .io_next_Q(bds_9_io_next_Q)
  );
  booth_div_substep bds_10 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_10_io_acc),
    .io_Q(bds_10_io_Q),
    .io_divisor(bds_10_io_divisor),
    .io_next_acc(bds_10_io_next_acc),
    .io_next_Q(bds_10_io_next_Q)
  );
  booth_div_substep bds_11 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_11_io_acc),
    .io_Q(bds_11_io_Q),
    .io_divisor(bds_11_io_divisor),
    .io_next_acc(bds_11_io_next_acc),
    .io_next_Q(bds_11_io_next_Q)
  );
  booth_div_substep bds_12 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_12_io_acc),
    .io_Q(bds_12_io_Q),
    .io_divisor(bds_12_io_divisor),
    .io_next_acc(bds_12_io_next_acc),
    .io_next_Q(bds_12_io_next_Q)
  );
  booth_div_substep bds_13 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_13_io_acc),
    .io_Q(bds_13_io_Q),
    .io_divisor(bds_13_io_divisor),
    .io_next_acc(bds_13_io_next_acc),
    .io_next_Q(bds_13_io_next_Q)
  );
  booth_div_substep bds_14 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_14_io_acc),
    .io_Q(bds_14_io_Q),
    .io_divisor(bds_14_io_divisor),
    .io_next_acc(bds_14_io_next_acc),
    .io_next_Q(bds_14_io_next_Q)
  );
  booth_div_substep bds_15 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_15_io_acc),
    .io_Q(bds_15_io_Q),
    .io_divisor(bds_15_io_divisor),
    .io_next_acc(bds_15_io_next_acc),
    .io_next_Q(bds_15_io_next_Q)
  );
  booth_div_substep bds_16 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_16_io_acc),
    .io_Q(bds_16_io_Q),
    .io_divisor(bds_16_io_divisor),
    .io_next_acc(bds_16_io_next_acc),
    .io_next_Q(bds_16_io_next_Q)
  );
  booth_div_substep bds_17 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_17_io_acc),
    .io_Q(bds_17_io_Q),
    .io_divisor(bds_17_io_divisor),
    .io_next_acc(bds_17_io_next_acc),
    .io_next_Q(bds_17_io_next_Q)
  );
  booth_div_substep bds_18 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_18_io_acc),
    .io_Q(bds_18_io_Q),
    .io_divisor(bds_18_io_divisor),
    .io_next_acc(bds_18_io_next_acc),
    .io_next_Q(bds_18_io_next_Q)
  );
  booth_div_substep bds_19 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_19_io_acc),
    .io_Q(bds_19_io_Q),
    .io_divisor(bds_19_io_divisor),
    .io_next_acc(bds_19_io_next_acc),
    .io_next_Q(bds_19_io_next_Q)
  );
  booth_div_substep bds_20 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_20_io_acc),
    .io_Q(bds_20_io_Q),
    .io_divisor(bds_20_io_divisor),
    .io_next_acc(bds_20_io_next_acc),
    .io_next_Q(bds_20_io_next_Q)
  );
  booth_div_substep bds_21 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_21_io_acc),
    .io_Q(bds_21_io_Q),
    .io_divisor(bds_21_io_divisor),
    .io_next_acc(bds_21_io_next_acc),
    .io_next_Q(bds_21_io_next_Q)
  );
  booth_div_substep bds_22 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_22_io_acc),
    .io_Q(bds_22_io_Q),
    .io_divisor(bds_22_io_divisor),
    .io_next_acc(bds_22_io_next_acc),
    .io_next_Q(bds_22_io_next_Q)
  );
  booth_div_substep bds_23 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_23_io_acc),
    .io_Q(bds_23_io_Q),
    .io_divisor(bds_23_io_divisor),
    .io_next_acc(bds_23_io_next_acc),
    .io_next_Q(bds_23_io_next_Q)
  );
  booth_div_substep bds_24 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_24_io_acc),
    .io_Q(bds_24_io_Q),
    .io_divisor(bds_24_io_divisor),
    .io_next_acc(bds_24_io_next_acc),
    .io_next_Q(bds_24_io_next_Q)
  );
  booth_div_substep bds_25 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_25_io_acc),
    .io_Q(bds_25_io_Q),
    .io_divisor(bds_25_io_divisor),
    .io_next_acc(bds_25_io_next_acc),
    .io_next_Q(bds_25_io_next_Q)
  );
  booth_div_substep bds_26 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_26_io_acc),
    .io_Q(bds_26_io_Q),
    .io_divisor(bds_26_io_divisor),
    .io_next_acc(bds_26_io_next_acc),
    .io_next_Q(bds_26_io_next_Q)
  );
  booth_div_substep bds_27 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_27_io_acc),
    .io_Q(bds_27_io_Q),
    .io_divisor(bds_27_io_divisor),
    .io_next_acc(bds_27_io_next_acc),
    .io_next_Q(bds_27_io_next_Q)
  );
  booth_div_substep bds_28 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_28_io_acc),
    .io_Q(bds_28_io_Q),
    .io_divisor(bds_28_io_divisor),
    .io_next_acc(bds_28_io_next_acc),
    .io_next_Q(bds_28_io_next_Q)
  );
  booth_div_substep bds_29 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_29_io_acc),
    .io_Q(bds_29_io_Q),
    .io_divisor(bds_29_io_divisor),
    .io_next_acc(bds_29_io_next_acc),
    .io_next_Q(bds_29_io_next_Q)
  );
  booth_div_substep bds_30 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_30_io_acc),
    .io_Q(bds_30_io_Q),
    .io_divisor(bds_30_io_divisor),
    .io_next_acc(bds_30_io_next_acc),
    .io_next_Q(bds_30_io_next_Q)
  );
  booth_div_substep bds_31 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_31_io_acc),
    .io_Q(bds_31_io_Q),
    .io_divisor(bds_31_io_divisor),
    .io_next_acc(bds_31_io_next_acc),
    .io_next_Q(bds_31_io_next_Q)
  );
  booth_div_substep bds_32 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_32_io_acc),
    .io_Q(bds_32_io_Q),
    .io_divisor(bds_32_io_divisor),
    .io_next_acc(bds_32_io_next_acc),
    .io_next_Q(bds_32_io_next_Q)
  );
  booth_div_substep bds_33 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_33_io_acc),
    .io_Q(bds_33_io_Q),
    .io_divisor(bds_33_io_divisor),
    .io_next_acc(bds_33_io_next_acc),
    .io_next_Q(bds_33_io_next_Q)
  );
  booth_div_substep bds_34 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_34_io_acc),
    .io_Q(bds_34_io_Q),
    .io_divisor(bds_34_io_divisor),
    .io_next_acc(bds_34_io_next_acc),
    .io_next_Q(bds_34_io_next_Q)
  );
  booth_div_substep bds_35 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_35_io_acc),
    .io_Q(bds_35_io_Q),
    .io_divisor(bds_35_io_divisor),
    .io_next_acc(bds_35_io_next_acc),
    .io_next_Q(bds_35_io_next_Q)
  );
  booth_div_substep bds_36 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_36_io_acc),
    .io_Q(bds_36_io_Q),
    .io_divisor(bds_36_io_divisor),
    .io_next_acc(bds_36_io_next_acc),
    .io_next_Q(bds_36_io_next_Q)
  );
  booth_div_substep bds_37 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_37_io_acc),
    .io_Q(bds_37_io_Q),
    .io_divisor(bds_37_io_divisor),
    .io_next_acc(bds_37_io_next_acc),
    .io_next_Q(bds_37_io_next_Q)
  );
  booth_div_substep bds_38 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_38_io_acc),
    .io_Q(bds_38_io_Q),
    .io_divisor(bds_38_io_divisor),
    .io_next_acc(bds_38_io_next_acc),
    .io_next_Q(bds_38_io_next_Q)
  );
  booth_div_substep bds_39 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_39_io_acc),
    .io_Q(bds_39_io_Q),
    .io_divisor(bds_39_io_divisor),
    .io_next_acc(bds_39_io_next_acc),
    .io_next_Q(bds_39_io_next_Q)
  );
  booth_div_substep bds_40 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_40_io_acc),
    .io_Q(bds_40_io_Q),
    .io_divisor(bds_40_io_divisor),
    .io_next_acc(bds_40_io_next_acc),
    .io_next_Q(bds_40_io_next_Q)
  );
  booth_div_substep bds_41 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_41_io_acc),
    .io_Q(bds_41_io_Q),
    .io_divisor(bds_41_io_divisor),
    .io_next_acc(bds_41_io_next_acc),
    .io_next_Q(bds_41_io_next_Q)
  );
  booth_div_substep bds_42 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_42_io_acc),
    .io_Q(bds_42_io_Q),
    .io_divisor(bds_42_io_divisor),
    .io_next_acc(bds_42_io_next_acc),
    .io_next_Q(bds_42_io_next_Q)
  );
  booth_div_substep bds_43 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_43_io_acc),
    .io_Q(bds_43_io_Q),
    .io_divisor(bds_43_io_divisor),
    .io_next_acc(bds_43_io_next_acc),
    .io_next_Q(bds_43_io_next_Q)
  );
  booth_div_substep bds_44 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_44_io_acc),
    .io_Q(bds_44_io_Q),
    .io_divisor(bds_44_io_divisor),
    .io_next_acc(bds_44_io_next_acc),
    .io_next_Q(bds_44_io_next_Q)
  );
  booth_div_substep bds_45 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_45_io_acc),
    .io_Q(bds_45_io_Q),
    .io_divisor(bds_45_io_divisor),
    .io_next_acc(bds_45_io_next_acc),
    .io_next_Q(bds_45_io_next_Q)
  );
  booth_div_substep bds_46 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_46_io_acc),
    .io_Q(bds_46_io_Q),
    .io_divisor(bds_46_io_divisor),
    .io_next_acc(bds_46_io_next_acc),
    .io_next_Q(bds_46_io_next_Q)
  );
  booth_div_substep bds_47 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_47_io_acc),
    .io_Q(bds_47_io_Q),
    .io_divisor(bds_47_io_divisor),
    .io_next_acc(bds_47_io_next_acc),
    .io_next_Q(bds_47_io_next_Q)
  );
  booth_div_substep bds_48 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_48_io_acc),
    .io_Q(bds_48_io_Q),
    .io_divisor(bds_48_io_divisor),
    .io_next_acc(bds_48_io_next_acc),
    .io_next_Q(bds_48_io_next_Q)
  );
  booth_div_substep bds_49 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_49_io_acc),
    .io_Q(bds_49_io_Q),
    .io_divisor(bds_49_io_divisor),
    .io_next_acc(bds_49_io_next_acc),
    .io_next_Q(bds_49_io_next_Q)
  );
  booth_div_substep bds_50 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_50_io_acc),
    .io_Q(bds_50_io_Q),
    .io_divisor(bds_50_io_divisor),
    .io_next_acc(bds_50_io_next_acc),
    .io_next_Q(bds_50_io_next_Q)
  );
  booth_div_substep bds_51 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_51_io_acc),
    .io_Q(bds_51_io_Q),
    .io_divisor(bds_51_io_divisor),
    .io_next_acc(bds_51_io_next_acc),
    .io_next_Q(bds_51_io_next_Q)
  );
  booth_div_substep bds_52 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_52_io_acc),
    .io_Q(bds_52_io_Q),
    .io_divisor(bds_52_io_divisor),
    .io_next_acc(bds_52_io_next_acc),
    .io_next_Q(bds_52_io_next_Q)
  );
  booth_div_substep bds_53 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_53_io_acc),
    .io_Q(bds_53_io_Q),
    .io_divisor(bds_53_io_divisor),
    .io_next_acc(bds_53_io_next_acc),
    .io_next_Q(bds_53_io_next_Q)
  );
  booth_div_substep bds_54 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_54_io_acc),
    .io_Q(bds_54_io_Q),
    .io_divisor(bds_54_io_divisor),
    .io_next_acc(bds_54_io_next_acc),
    .io_next_Q(bds_54_io_next_Q)
  );
  booth_div_substep bds_55 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_55_io_acc),
    .io_Q(bds_55_io_Q),
    .io_divisor(bds_55_io_divisor),
    .io_next_acc(bds_55_io_next_acc),
    .io_next_Q(bds_55_io_next_Q)
  );
  booth_div_substep bds_56 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_56_io_acc),
    .io_Q(bds_56_io_Q),
    .io_divisor(bds_56_io_divisor),
    .io_next_acc(bds_56_io_next_acc),
    .io_next_Q(bds_56_io_next_Q)
  );
  booth_div_substep bds_57 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_57_io_acc),
    .io_Q(bds_57_io_Q),
    .io_divisor(bds_57_io_divisor),
    .io_next_acc(bds_57_io_next_acc),
    .io_next_Q(bds_57_io_next_Q)
  );
  booth_div_substep bds_58 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_58_io_acc),
    .io_Q(bds_58_io_Q),
    .io_divisor(bds_58_io_divisor),
    .io_next_acc(bds_58_io_next_acc),
    .io_next_Q(bds_58_io_next_Q)
  );
  booth_div_substep bds_59 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_59_io_acc),
    .io_Q(bds_59_io_Q),
    .io_divisor(bds_59_io_divisor),
    .io_next_acc(bds_59_io_next_acc),
    .io_next_Q(bds_59_io_next_Q)
  );
  booth_div_substep bds_60 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_60_io_acc),
    .io_Q(bds_60_io_Q),
    .io_divisor(bds_60_io_divisor),
    .io_next_acc(bds_60_io_next_acc),
    .io_next_Q(bds_60_io_next_Q)
  );
  booth_div_substep bds_61 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_61_io_acc),
    .io_Q(bds_61_io_Q),
    .io_divisor(bds_61_io_divisor),
    .io_next_acc(bds_61_io_next_acc),
    .io_next_Q(bds_61_io_next_Q)
  );
  booth_div_substep bds_62 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_62_io_acc),
    .io_Q(bds_62_io_Q),
    .io_divisor(bds_62_io_divisor),
    .io_next_acc(bds_62_io_next_acc),
    .io_next_Q(bds_62_io_next_Q)
  );
  booth_div_substep bds_63 ( // @[booth_divider.scala 51:33]
    .io_acc(bds_63_io_acc),
    .io_Q(bds_63_io_Q),
    .io_divisor(bds_63_io_divisor),
    .io_next_acc(bds_63_io_next_acc),
    .io_next_Q(bds_63_io_next_Q)
  );
  assign io_quotient = neg_quotient ? _T_26 : quotientTemp; // @[booth_divider.scala 69:83]
  assign io_remainder = _T_16 ? _T_35 : remainderTemp; // @[booth_divider.scala 70:112]
  assign bds_0_io_acc = 64'h0; // @[booth_divider.scala 43:19 booth_divider.scala 49:13]
  assign bds_0_io_Q = io_signed & io_dividend[63] ? dividend_comp : io_dividend; // @[booth_divider.scala 29:56 booth_divider.scala 30:21 booth_divider.scala 32:21]
  assign bds_0_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_1_io_acc = bds_0_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_1_io_Q = bds_0_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_1_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_2_io_acc = bds_1_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_2_io_Q = bds_1_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_2_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_3_io_acc = bds_2_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_3_io_Q = bds_2_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_3_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_4_io_acc = bds_3_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_4_io_Q = bds_3_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_4_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_5_io_acc = bds_4_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_5_io_Q = bds_4_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_5_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_6_io_acc = bds_5_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_6_io_Q = bds_5_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_6_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_7_io_acc = bds_6_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_7_io_Q = bds_6_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_7_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_8_io_acc = bds_7_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_8_io_Q = bds_7_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_8_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_9_io_acc = bds_8_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_9_io_Q = bds_8_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_9_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_10_io_acc = bds_9_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_10_io_Q = bds_9_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_10_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_11_io_acc = bds_10_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_11_io_Q = bds_10_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_11_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_12_io_acc = bds_11_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_12_io_Q = bds_11_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_12_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_13_io_acc = bds_12_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_13_io_Q = bds_12_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_13_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_14_io_acc = bds_13_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_14_io_Q = bds_13_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_14_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_15_io_acc = bds_14_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_15_io_Q = bds_14_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_15_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_16_io_acc = bds_15_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_16_io_Q = bds_15_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_16_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_17_io_acc = bds_16_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_17_io_Q = bds_16_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_17_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_18_io_acc = bds_17_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_18_io_Q = bds_17_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_18_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_19_io_acc = bds_18_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_19_io_Q = bds_18_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_19_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_20_io_acc = bds_19_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_20_io_Q = bds_19_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_20_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_21_io_acc = bds_20_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_21_io_Q = bds_20_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_21_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_22_io_acc = bds_21_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_22_io_Q = bds_21_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_22_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_23_io_acc = bds_22_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_23_io_Q = bds_22_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_23_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_24_io_acc = bds_23_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_24_io_Q = bds_23_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_24_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_25_io_acc = bds_24_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_25_io_Q = bds_24_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_25_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_26_io_acc = bds_25_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_26_io_Q = bds_25_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_26_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_27_io_acc = bds_26_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_27_io_Q = bds_26_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_27_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_28_io_acc = bds_27_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_28_io_Q = bds_27_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_28_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_29_io_acc = bds_28_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_29_io_Q = bds_28_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_29_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_30_io_acc = bds_29_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_30_io_Q = bds_29_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_30_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_31_io_acc = bds_30_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_31_io_Q = bds_30_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_31_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_32_io_acc = bds_31_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_32_io_Q = bds_31_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_32_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_33_io_acc = bds_32_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_33_io_Q = bds_32_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_33_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_34_io_acc = bds_33_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_34_io_Q = bds_33_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_34_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_35_io_acc = bds_34_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_35_io_Q = bds_34_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_35_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_36_io_acc = bds_35_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_36_io_Q = bds_35_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_36_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_37_io_acc = bds_36_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_37_io_Q = bds_36_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_37_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_38_io_acc = bds_37_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_38_io_Q = bds_37_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_38_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_39_io_acc = bds_38_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_39_io_Q = bds_38_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_39_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_40_io_acc = bds_39_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_40_io_Q = bds_39_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_40_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_41_io_acc = bds_40_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_41_io_Q = bds_40_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_41_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_42_io_acc = bds_41_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_42_io_Q = bds_41_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_42_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_43_io_acc = bds_42_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_43_io_Q = bds_42_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_43_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_44_io_acc = bds_43_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_44_io_Q = bds_43_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_44_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_45_io_acc = bds_44_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_45_io_Q = bds_44_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_45_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_46_io_acc = bds_45_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_46_io_Q = bds_45_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_46_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_47_io_acc = bds_46_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_47_io_Q = bds_46_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_47_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_48_io_acc = bds_47_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_48_io_Q = bds_47_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_48_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_49_io_acc = bds_48_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_49_io_Q = bds_48_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_49_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_50_io_acc = bds_49_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_50_io_Q = bds_49_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_50_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_51_io_acc = bds_50_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_51_io_Q = bds_50_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_51_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_52_io_acc = bds_51_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_52_io_Q = bds_51_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_52_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_53_io_acc = bds_52_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_53_io_Q = bds_52_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_53_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_54_io_acc = bds_53_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_54_io_Q = bds_53_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_54_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_55_io_acc = bds_54_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_55_io_Q = bds_54_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_55_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_56_io_acc = bds_55_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_56_io_Q = bds_55_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_56_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_57_io_acc = bds_56_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_57_io_Q = bds_56_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_57_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_58_io_acc = bds_57_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_58_io_Q = bds_57_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_58_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_59_io_acc = bds_58_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_59_io_Q = bds_58_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_59_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_60_io_acc = bds_59_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_60_io_Q = bds_59_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_60_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_61_io_acc = bds_60_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_61_io_Q = bds_60_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_61_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_62_io_acc = bds_61_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_62_io_Q = bds_61_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_62_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
  assign bds_63_io_acc = bds_62_io_next_acc; // @[booth_divider.scala 43:19 booth_divider.scala 57:29]
  assign bds_63_io_Q = bds_62_io_next_Q; // @[booth_divider.scala 42:17 booth_divider.scala 58:29]
  assign bds_63_io_divisor = io_signed & io_divisor[63] ? divisor_comp : io_divisor; // @[booth_divider.scala 35:55 booth_divider.scala 36:20 booth_divider.scala 38:20]
endmodule
